module cam_allocator_neo(
  input         clock,
  input         reset,
  output [1:0]  io_res_search_out,
  input         io_res_search_en,
  output [11:0] io_res_search_out_start_0,
  output [11:0] io_res_search_out_start_1,
  input  [12:0] io_res_search_size,
  input         io_cam_wr_en,
  input  [1:0]  io_cam_wr_addr,
  input  [12:0] io_cam_wr_data,
  input  [11:0] io_cam_wr_start
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  res_search_en_i; // @[cam_allocator_neo.scala 17:34]
  reg [12:0] res_search_size_i; // @[cam_allocator_neo.scala 18:36]
  reg  cam_valid_entry_0; // @[cam_allocator_neo.scala 19:34]
  reg  cam_valid_entry_1; // @[cam_allocator_neo.scala 19:34]
  reg [12:0] cam_ram_0; // @[cam_allocator_neo.scala 20:26]
  reg [12:0] cam_ram_1; // @[cam_allocator_neo.scala 20:26]
  reg [11:0] cam_ram_start_0; // @[cam_allocator_neo.scala 21:32]
  reg [11:0] cam_ram_start_1; // @[cam_allocator_neo.scala 21:32]
  wire  _T_2 = cam_ram_0 >= res_search_size_i; // @[cam_allocator_neo.scala 37:33]
  wire  _GEN_1 = ~cam_valid_entry_0 | _T_2; // @[cam_allocator_neo.scala 33:38 34:35]
  wire  decoded_output_0 = ~res_search_en_i ? 1'h0 : _GEN_1; // @[cam_allocator_neo.scala 29:31 30:31]
  wire  _T_5 = cam_ram_1 >= res_search_size_i; // @[cam_allocator_neo.scala 37:33]
  wire  _GEN_4 = ~cam_valid_entry_1 | _T_5; // @[cam_allocator_neo.scala 33:38 34:35]
  wire  decoded_output_1 = ~res_search_en_i ? 1'h0 : _GEN_4; // @[cam_allocator_neo.scala 29:31 30:31]
  wire  _GEN_10 = ~io_cam_wr_addr[0] | cam_valid_entry_0; // @[cam_allocator_neo.scala 19:34 52:{41,41}]
  wire  _GEN_11 = io_cam_wr_addr[0] | cam_valid_entry_1; // @[cam_allocator_neo.scala 19:34 52:{41,41}]
  assign io_res_search_out = {decoded_output_1,decoded_output_0}; // @[cam_allocator_neo.scala 54:41]
  assign io_res_search_out_start_0 = cam_ram_start_0; // @[cam_allocator_neo.scala 23:38]
  assign io_res_search_out_start_1 = cam_ram_start_1; // @[cam_allocator_neo.scala 23:38]
  always @(posedge clock) begin
    if (reset) begin // @[cam_allocator_neo.scala 17:34]
      res_search_en_i <= 1'h0; // @[cam_allocator_neo.scala 17:34]
    end else begin
      res_search_en_i <= io_res_search_en; // @[cam_allocator_neo.scala 26:21]
    end
    if (reset) begin // @[cam_allocator_neo.scala 18:36]
      res_search_size_i <= 13'h0; // @[cam_allocator_neo.scala 18:36]
    end else begin
      res_search_size_i <= io_res_search_size; // @[cam_allocator_neo.scala 27:23]
    end
    if (reset) begin // @[cam_allocator_neo.scala 19:34]
      cam_valid_entry_0 <= 1'h0; // @[cam_allocator_neo.scala 19:34]
    end else if (io_cam_wr_en) begin // @[cam_allocator_neo.scala 48:23]
      cam_valid_entry_0 <= _GEN_10;
    end
    if (reset) begin // @[cam_allocator_neo.scala 19:34]
      cam_valid_entry_1 <= 1'h0; // @[cam_allocator_neo.scala 19:34]
    end else if (io_cam_wr_en) begin // @[cam_allocator_neo.scala 48:23]
      cam_valid_entry_1 <= _GEN_11;
    end
    if (reset) begin // @[cam_allocator_neo.scala 20:26]
      cam_ram_0 <= 13'h0; // @[cam_allocator_neo.scala 20:26]
    end else if (io_cam_wr_en) begin // @[cam_allocator_neo.scala 48:23]
      if (~io_cam_wr_addr[0]) begin // @[cam_allocator_neo.scala 50:33]
        cam_ram_0 <= io_cam_wr_data; // @[cam_allocator_neo.scala 50:33]
      end
    end
    if (reset) begin // @[cam_allocator_neo.scala 20:26]
      cam_ram_1 <= 13'h0; // @[cam_allocator_neo.scala 20:26]
    end else if (io_cam_wr_en) begin // @[cam_allocator_neo.scala 48:23]
      if (io_cam_wr_addr[0]) begin // @[cam_allocator_neo.scala 50:33]
        cam_ram_1 <= io_cam_wr_data; // @[cam_allocator_neo.scala 50:33]
      end
    end
    if (reset) begin // @[cam_allocator_neo.scala 21:32]
      cam_ram_start_0 <= 12'h0; // @[cam_allocator_neo.scala 21:32]
    end else if (io_cam_wr_en) begin // @[cam_allocator_neo.scala 48:23]
      if (~io_cam_wr_addr[0]) begin // @[cam_allocator_neo.scala 51:39]
        cam_ram_start_0 <= io_cam_wr_start; // @[cam_allocator_neo.scala 51:39]
      end
    end
    if (reset) begin // @[cam_allocator_neo.scala 21:32]
      cam_ram_start_1 <= 12'h0; // @[cam_allocator_neo.scala 21:32]
    end else if (io_cam_wr_en) begin // @[cam_allocator_neo.scala 48:23]
      if (io_cam_wr_addr[0]) begin // @[cam_allocator_neo.scala 51:39]
        cam_ram_start_1 <= io_cam_wr_start; // @[cam_allocator_neo.scala 51:39]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  res_search_en_i = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  res_search_size_i = _RAND_1[12:0];
  _RAND_2 = {1{`RANDOM}};
  cam_valid_entry_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cam_valid_entry_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cam_ram_0 = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  cam_ram_1 = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  cam_ram_start_0 = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  cam_ram_start_1 = _RAND_7[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cam_allocator(
  input        clock,
  input        reset,
  output [1:0] io_res_search_out,
  input        io_res_search_en,
  input  [3:0] io_res_search_size,
  input        io_cam_wr_en,
  input  [1:0] io_cam_wr_addr,
  input  [3:0] io_cam_wr_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  res_search_en_i; // @[cam_allocator.scala 16:34]
  reg [3:0] res_search_size_i; // @[cam_allocator.scala 17:36]
  reg  cam_valid_entry_0; // @[cam_allocator.scala 18:34]
  reg  cam_valid_entry_1; // @[cam_allocator.scala 18:34]
  reg [3:0] cam_ram_0; // @[cam_allocator.scala 19:26]
  reg [3:0] cam_ram_1; // @[cam_allocator.scala 19:26]
  wire  _T_2 = cam_ram_0 >= res_search_size_i; // @[cam_allocator.scala 32:33]
  wire  _GEN_1 = ~cam_valid_entry_0 | _T_2; // @[cam_allocator.scala 28:38 29:35]
  wire  decoded_output_0 = ~res_search_en_i ? 1'h0 : _GEN_1; // @[cam_allocator.scala 24:31 25:31]
  wire  _T_5 = cam_ram_1 >= res_search_size_i; // @[cam_allocator.scala 32:33]
  wire  _GEN_4 = ~cam_valid_entry_1 | _T_5; // @[cam_allocator.scala 28:38 29:35]
  wire  decoded_output_1 = ~res_search_en_i ? 1'h0 : _GEN_4; // @[cam_allocator.scala 24:31 25:31]
  wire  _GEN_8 = ~io_cam_wr_addr[0] | cam_valid_entry_0; // @[cam_allocator.scala 18:34 43:{41,41}]
  wire  _GEN_9 = io_cam_wr_addr[0] | cam_valid_entry_1; // @[cam_allocator.scala 18:34 43:{41,41}]
  assign io_res_search_out = {decoded_output_1,decoded_output_0}; // @[cam_allocator.scala 45:41]
  always @(posedge clock) begin
    if (reset) begin // @[cam_allocator.scala 16:34]
      res_search_en_i <= 1'h0; // @[cam_allocator.scala 16:34]
    end else begin
      res_search_en_i <= io_res_search_en; // @[cam_allocator.scala 21:21]
    end
    if (reset) begin // @[cam_allocator.scala 17:36]
      res_search_size_i <= 4'h0; // @[cam_allocator.scala 17:36]
    end else begin
      res_search_size_i <= io_res_search_size; // @[cam_allocator.scala 22:23]
    end
    if (reset) begin // @[cam_allocator.scala 18:34]
      cam_valid_entry_0 <= 1'h0; // @[cam_allocator.scala 18:34]
    end else if (io_cam_wr_en) begin // @[cam_allocator.scala 41:23]
      cam_valid_entry_0 <= _GEN_8;
    end
    if (reset) begin // @[cam_allocator.scala 18:34]
      cam_valid_entry_1 <= 1'h0; // @[cam_allocator.scala 18:34]
    end else if (io_cam_wr_en) begin // @[cam_allocator.scala 41:23]
      cam_valid_entry_1 <= _GEN_9;
    end
    if (reset) begin // @[cam_allocator.scala 19:26]
      cam_ram_0 <= 4'h0; // @[cam_allocator.scala 19:26]
    end else if (io_cam_wr_en) begin // @[cam_allocator.scala 41:23]
      if (~io_cam_wr_addr[0]) begin // @[cam_allocator.scala 42:33]
        cam_ram_0 <= io_cam_wr_data; // @[cam_allocator.scala 42:33]
      end
    end
    if (reset) begin // @[cam_allocator.scala 19:26]
      cam_ram_1 <= 4'h0; // @[cam_allocator.scala 19:26]
    end else if (io_cam_wr_en) begin // @[cam_allocator.scala 41:23]
      if (io_cam_wr_addr[0]) begin // @[cam_allocator.scala 42:33]
        cam_ram_1 <= io_cam_wr_data; // @[cam_allocator.scala 42:33]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  res_search_en_i = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  res_search_size_i = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  cam_valid_entry_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cam_valid_entry_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cam_ram_0 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  cam_ram_1 = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module prefer_select(
  input        io_signal_0,
  input        io_signal_1,
  input  [1:0] io_prefer,
  output       io_valid,
  output [1:0] io_id
);
  wire [2:0] _GEN_20 = {{1'd0}, io_prefer}; // @[prefer_select.scala 17:36]
  wire [2:0] _T_1 = 3'h1 + _GEN_20; // @[prefer_select.scala 17:36]
  wire [2:0] _T_6 = _T_1 - 3'h2; // @[prefer_select.scala 18:62]
  wire  _GEN_1 = _T_6[0] ? io_signal_1 : io_signal_0; // @[prefer_select.scala 18:{91,91}]
  wire [2:0] _GEN_3 = _GEN_1 ? _T_6 : 3'h0; // @[prefer_select.scala 15:14 18:91 20:26]
  wire [1:0] _T_9 = 2'h1 + io_prefer; // @[prefer_select.scala 24:32]
  wire  _GEN_5 = _T_9[0] ? io_signal_1 : io_signal_0; // @[prefer_select.scala 24:{45,45}]
  wire [1:0] _GEN_7 = _GEN_5 ? _T_9 : 2'h0; // @[prefer_select.scala 15:14 24:45 26:26]
  wire  _GEN_8 = _T_1 >= 3'h2 ? _GEN_1 : _GEN_5; // @[prefer_select.scala 17:77]
  wire [2:0] _GEN_9 = _T_1 >= 3'h2 ? _GEN_3 : {{1'd0}, _GEN_7}; // @[prefer_select.scala 17:77]
  wire [2:0] _T_12 = 3'h2 + _GEN_20; // @[prefer_select.scala 17:36]
  wire [2:0] _T_17 = _T_12 - 3'h2; // @[prefer_select.scala 18:62]
  wire  _GEN_11 = _T_17[0] ? io_signal_1 : io_signal_0; // @[prefer_select.scala 18:{91,91}]
  wire  _GEN_12 = _GEN_11 | _GEN_8; // @[prefer_select.scala 18:91 19:23]
  wire [2:0] _GEN_13 = _GEN_11 ? _T_17 : _GEN_9; // @[prefer_select.scala 18:91 20:26]
  wire [1:0] _T_20 = 2'h2 + io_prefer; // @[prefer_select.scala 24:32]
  wire  _GEN_15 = _T_20[0] ? io_signal_1 : io_signal_0; // @[prefer_select.scala 24:{45,45}]
  wire  _GEN_16 = _GEN_15 | _GEN_8; // @[prefer_select.scala 24:45 25:23]
  wire [2:0] _GEN_17 = _GEN_15 ? {{1'd0}, _T_20} : _GEN_9; // @[prefer_select.scala 24:45 26:26]
  wire [2:0] found_id = _T_12 >= 3'h2 ? _GEN_13 : _GEN_17; // @[prefer_select.scala 17:77]
  assign io_valid = _T_12 >= 3'h2 ? _GEN_12 : _GEN_16; // @[prefer_select.scala 17:77]
  assign io_id = found_id[1:0]; // @[prefer_select.scala 31:22]
endmodule
module allocator_neo(
  input         clock,
  input         reset,
  output        io_allocator_cu_valid,
  output        io_allocator_cu_rejected,
  output [4:0]  io_allocator_wg_id_out,
  output [1:0]  io_allocator_cu_id_out,
  output [2:0]  io_allocator_wf_count,
  output [12:0] io_allocator_vgpr_size_out,
  output [12:0] io_allocator_sgpr_size_out,
  output [12:0] io_allocator_lds_size_out,
  output [11:0] io_allocator_vgpr_start_out,
  output [11:0] io_allocator_sgpr_start_out,
  output [11:0] io_allocator_lds_start_out,
  input  [4:0]  io_inflight_wg_buffer_alloc_wg_id,
  input  [2:0]  io_inflight_wg_buffer_alloc_num_wf,
  input  [12:0] io_inflight_wg_buffer_alloc_vgpr_size,
  input  [12:0] io_inflight_wg_buffer_alloc_sgpr_size,
  input  [12:0] io_inflight_wg_buffer_alloc_lds_size,
  input  [1:0]  io_dis_controller_cu_busy,
  input         io_dis_controller_alloc_ack,
  input         io_dis_controller_start_alloc,
  input         io_grt_cam_up_valid,
  input  [1:0]  io_grt_cam_up_cu_id,
  input  [11:0] io_grt_cam_up_vgpr_strt,
  input  [12:0] io_grt_cam_up_vgpr_size,
  input  [11:0] io_grt_cam_up_sgpr_strt,
  input  [12:0] io_grt_cam_up_sgpr_size,
  input  [11:0] io_grt_cam_up_lds_strt,
  input  [12:0] io_grt_cam_up_lds_size,
  input  [2:0]  io_grt_cam_up_wf_count,
  input  [2:0]  io_grt_cam_up_wg_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
`endif // RANDOMIZE_REG_INIT
  wire  vgpr_cam_clock; // @[allocator_neo.scala 129:26]
  wire  vgpr_cam_reset; // @[allocator_neo.scala 129:26]
  wire [1:0] vgpr_cam_io_res_search_out; // @[allocator_neo.scala 129:26]
  wire  vgpr_cam_io_res_search_en; // @[allocator_neo.scala 129:26]
  wire [11:0] vgpr_cam_io_res_search_out_start_0; // @[allocator_neo.scala 129:26]
  wire [11:0] vgpr_cam_io_res_search_out_start_1; // @[allocator_neo.scala 129:26]
  wire [12:0] vgpr_cam_io_res_search_size; // @[allocator_neo.scala 129:26]
  wire  vgpr_cam_io_cam_wr_en; // @[allocator_neo.scala 129:26]
  wire [1:0] vgpr_cam_io_cam_wr_addr; // @[allocator_neo.scala 129:26]
  wire [12:0] vgpr_cam_io_cam_wr_data; // @[allocator_neo.scala 129:26]
  wire [11:0] vgpr_cam_io_cam_wr_start; // @[allocator_neo.scala 129:26]
  wire  sgpr_cam_clock; // @[allocator_neo.scala 130:26]
  wire  sgpr_cam_reset; // @[allocator_neo.scala 130:26]
  wire [1:0] sgpr_cam_io_res_search_out; // @[allocator_neo.scala 130:26]
  wire  sgpr_cam_io_res_search_en; // @[allocator_neo.scala 130:26]
  wire [11:0] sgpr_cam_io_res_search_out_start_0; // @[allocator_neo.scala 130:26]
  wire [11:0] sgpr_cam_io_res_search_out_start_1; // @[allocator_neo.scala 130:26]
  wire [12:0] sgpr_cam_io_res_search_size; // @[allocator_neo.scala 130:26]
  wire  sgpr_cam_io_cam_wr_en; // @[allocator_neo.scala 130:26]
  wire [1:0] sgpr_cam_io_cam_wr_addr; // @[allocator_neo.scala 130:26]
  wire [12:0] sgpr_cam_io_cam_wr_data; // @[allocator_neo.scala 130:26]
  wire [11:0] sgpr_cam_io_cam_wr_start; // @[allocator_neo.scala 130:26]
  wire  lds_cam_clock; // @[allocator_neo.scala 131:25]
  wire  lds_cam_reset; // @[allocator_neo.scala 131:25]
  wire [1:0] lds_cam_io_res_search_out; // @[allocator_neo.scala 131:25]
  wire  lds_cam_io_res_search_en; // @[allocator_neo.scala 131:25]
  wire [11:0] lds_cam_io_res_search_out_start_0; // @[allocator_neo.scala 131:25]
  wire [11:0] lds_cam_io_res_search_out_start_1; // @[allocator_neo.scala 131:25]
  wire [12:0] lds_cam_io_res_search_size; // @[allocator_neo.scala 131:25]
  wire  lds_cam_io_cam_wr_en; // @[allocator_neo.scala 131:25]
  wire [1:0] lds_cam_io_cam_wr_addr; // @[allocator_neo.scala 131:25]
  wire [12:0] lds_cam_io_cam_wr_data; // @[allocator_neo.scala 131:25]
  wire [11:0] lds_cam_io_cam_wr_start; // @[allocator_neo.scala 131:25]
  wire  wf_cam_clock; // @[allocator_neo.scala 132:24]
  wire  wf_cam_reset; // @[allocator_neo.scala 132:24]
  wire [1:0] wf_cam_io_res_search_out; // @[allocator_neo.scala 132:24]
  wire  wf_cam_io_res_search_en; // @[allocator_neo.scala 132:24]
  wire [3:0] wf_cam_io_res_search_size; // @[allocator_neo.scala 132:24]
  wire  wf_cam_io_cam_wr_en; // @[allocator_neo.scala 132:24]
  wire [1:0] wf_cam_io_cam_wr_addr; // @[allocator_neo.scala 132:24]
  wire [3:0] wf_cam_io_cam_wr_data; // @[allocator_neo.scala 132:24]
  wire  wg_cam_clock; // @[allocator_neo.scala 133:24]
  wire  wg_cam_reset; // @[allocator_neo.scala 133:24]
  wire [1:0] wg_cam_io_res_search_out; // @[allocator_neo.scala 133:24]
  wire  wg_cam_io_res_search_en; // @[allocator_neo.scala 133:24]
  wire [3:0] wg_cam_io_res_search_size; // @[allocator_neo.scala 133:24]
  wire  wg_cam_io_cam_wr_en; // @[allocator_neo.scala 133:24]
  wire [1:0] wg_cam_io_cam_wr_addr; // @[allocator_neo.scala 133:24]
  wire [3:0] wg_cam_io_cam_wr_data; // @[allocator_neo.scala 133:24]
  wire  prefer_select_io_signal_0; // @[allocator_neo.scala 303:31]
  wire  prefer_select_io_signal_1; // @[allocator_neo.scala 303:31]
  wire [1:0] prefer_select_io_prefer; // @[allocator_neo.scala 303:31]
  wire  prefer_select_io_valid; // @[allocator_neo.scala 303:31]
  wire [1:0] prefer_select_io_id; // @[allocator_neo.scala 303:31]
  reg  alloc_valid_i; // @[allocator_neo.scala 42:32]
  reg [4:0] alloc_wg_id_i; // @[allocator_neo.scala 43:32]
  reg [2:0] alloc_num_wf_i; // @[allocator_neo.scala 44:33]
  reg [12:0] alloc_vgpr_size_i; // @[allocator_neo.scala 45:36]
  reg [12:0] alloc_sgpr_size_i; // @[allocator_neo.scala 46:36]
  reg [12:0] alloc_lds_size_i; // @[allocator_neo.scala 47:35]
  reg [1:0] dis_controller_cu_busy_i; // @[allocator_neo.scala 48:43]
  reg  cam_up_valid_i; // @[allocator_neo.scala 50:33]
  reg [1:0] cam_up_cu_id_i; // @[allocator_neo.scala 51:33]
  reg [11:0] cam_up_vgpr_strt_i; // @[allocator_neo.scala 52:37]
  reg [12:0] cam_up_vgpr_size_i; // @[allocator_neo.scala 53:37]
  reg [11:0] cam_up_sgpr_strt_i; // @[allocator_neo.scala 54:37]
  reg [12:0] cam_up_sgpr_size_i; // @[allocator_neo.scala 55:37]
  reg [11:0] cam_up_lds_strt_i; // @[allocator_neo.scala 56:36]
  reg [12:0] cam_up_lds_size_i; // @[allocator_neo.scala 57:36]
  reg [2:0] cam_up_wf_count_i; // @[allocator_neo.scala 58:36]
  reg [2:0] cam_up_wg_count_i; // @[allocator_neo.scala 59:36]
  reg  cam_wait_valid; // @[allocator_neo.scala 70:33]
  reg [4:0] cam_wait_wg_id; // @[allocator_neo.scala 71:33]
  reg [2:0] cam_wait_wf_count; // @[allocator_neo.scala 72:36]
  reg [12:0] cam_wait_vgpr_size; // @[allocator_neo.scala 73:37]
  reg [12:0] cam_wait_sgpr_size; // @[allocator_neo.scala 74:37]
  reg [12:0] cam_wait_lds_size; // @[allocator_neo.scala 75:36]
  reg [1:0] cam_wait_dis_controller_cu_busy; // @[allocator_neo.scala 76:50]
  reg  anded_cam_out_valid; // @[allocator_neo.scala 79:38]
  reg [1:0] anded_cam_out; // @[allocator_neo.scala 80:32]
  reg [4:0] anded_cam_wg_id; // @[allocator_neo.scala 81:34]
  reg [2:0] anded_cam_wf_count; // @[allocator_neo.scala 82:37]
  reg [12:0] anded_cam_vgpr_size; // @[allocator_neo.scala 83:38]
  reg [12:0] anded_cam_sgpr_size; // @[allocator_neo.scala 84:38]
  reg [12:0] anded_cam_lds_size; // @[allocator_neo.scala 85:37]
  reg  encoded_cu_out_valid; // @[allocator_neo.scala 88:39]
  reg  encoded_cu_found_valid; // @[allocator_neo.scala 89:41]
  reg [1:0] encoded_cu_id; // @[allocator_neo.scala 91:32]
  reg [4:0] encoded_cu_wg_id; // @[allocator_neo.scala 93:35]
  reg [2:0] encoded_wf_count; // @[allocator_neo.scala 94:35]
  reg [12:0] encoded_vgpr_size; // @[allocator_neo.scala 95:36]
  reg [12:0] encoded_sgpr_size; // @[allocator_neo.scala 96:36]
  reg [12:0] encoded_lds_size; // @[allocator_neo.scala 97:35]
  reg [11:0] encoded_vgpr_start; // @[allocator_neo.scala 98:37]
  reg [11:0] encoded_sgpr_start; // @[allocator_neo.scala 99:37]
  reg [11:0] encoded_lds_start; // @[allocator_neo.scala 100:36]
  reg  size_ram_valid; // @[allocator_neo.scala 103:33]
  reg  size_ram_cu_id_found; // @[allocator_neo.scala 104:39]
  reg [1:0] cu_id_out; // @[allocator_neo.scala 105:28]
  reg [11:0] vgpr_start_out; // @[allocator_neo.scala 106:33]
  reg [11:0] sgpr_start_out; // @[allocator_neo.scala 107:33]
  reg [11:0] lds_start_out; // @[allocator_neo.scala 108:32]
  reg [4:0] wg_id_out; // @[allocator_neo.scala 109:28]
  reg [2:0] wf_count_out; // @[allocator_neo.scala 110:31]
  reg [12:0] vgpr_size_out; // @[allocator_neo.scala 111:32]
  reg [12:0] sgpr_size_out; // @[allocator_neo.scala 112:32]
  reg [12:0] lds_size_out; // @[allocator_neo.scala 113:31]
  reg  cu_initialized_0; // @[allocator_neo.scala 125:33]
  reg  cu_initialized_1; // @[allocator_neo.scala 125:33]
  reg  pipeline_waiting; // @[allocator_neo.scala 127:35]
  wire  _T = ~pipeline_waiting; // @[allocator_neo.scala 193:36]
  wire  _GEN_0 = encoded_cu_found_valid & ~pipeline_waiting | pipeline_waiting; // @[allocator_neo.scala 193:54 194:26 127:35]
  wire [1:0] vgpr_search_out = vgpr_cam_io_res_search_out; // @[allocator_neo.scala 141:21 63:31]
  wire [1:0] sgpr_search_out = sgpr_cam_io_res_search_out; // @[allocator_neo.scala 152:21 64:31]
  wire [1:0] _anded_cam_out_T = vgpr_search_out & sgpr_search_out; // @[allocator_neo.scala 221:42]
  wire [1:0] lds_search_out = lds_cam_io_res_search_out; // @[allocator_neo.scala 163:20 65:30]
  wire [1:0] _anded_cam_out_T_1 = _anded_cam_out_T & lds_search_out; // @[allocator_neo.scala 221:60]
  wire [1:0] wf_search_out = wf_cam_io_res_search_out; // @[allocator_neo.scala 175:19 66:29]
  wire [1:0] _anded_cam_out_T_2 = _anded_cam_out_T_1 & wf_search_out; // @[allocator_neo.scala 221:77]
  wire [1:0] wg_search_out = wg_cam_io_res_search_out; // @[allocator_neo.scala 183:19 67:29]
  wire [1:0] _anded_cam_out_T_3 = _anded_cam_out_T_2 & wg_search_out; // @[allocator_neo.scala 221:93]
  wire [1:0] _anded_cam_out_T_4 = ~cam_wait_dis_controller_cu_busy; // @[allocator_neo.scala 221:111]
  wire [1:0] _anded_cam_out_T_5 = _anded_cam_out_T_3 & _anded_cam_out_T_4; // @[allocator_neo.scala 221:109]
  wire  encoded_cu_found_valid_comb = prefer_select_io_valid; // @[allocator_neo.scala 310:33 90:43]
  wire [1:0] encoded_cu_id_comb = prefer_select_io_id; // @[allocator_neo.scala 311:24 92:34]
  wire [11:0] lds_cam_start_vec_1 = lds_cam_io_res_search_out_start_1; // @[allocator_neo.scala 136:33 164:23]
  wire [11:0] lds_cam_start_vec_0 = lds_cam_io_res_search_out_start_0; // @[allocator_neo.scala 136:33 164:23]
  wire [11:0] vgpr_cam_start_vec_1 = vgpr_cam_io_res_search_out_start_1; // @[allocator_neo.scala 134:34 142:24]
  wire [11:0] vgpr_cam_start_vec_0 = vgpr_cam_io_res_search_out_start_0; // @[allocator_neo.scala 134:34 142:24]
  wire [11:0] sgpr_cam_start_vec_1 = sgpr_cam_io_res_search_out_start_1; // @[allocator_neo.scala 135:34 153:24]
  wire [11:0] sgpr_cam_start_vec_0 = sgpr_cam_io_res_search_out_start_0; // @[allocator_neo.scala 135:34 153:24]
  wire  _GEN_45 = ~cam_up_cu_id_i[0] | cu_initialized_0; // @[allocator_neo.scala 125:33 264:{40,40}]
  wire  _GEN_46 = cam_up_cu_id_i[0] | cu_initialized_1; // @[allocator_neo.scala 125:33 264:{40,40}]
  wire  _GEN_50 = cu_id_out[0] ? cu_initialized_1 : cu_initialized_0; // @[allocator_neo.scala 280:{10,10}]
  cam_allocator_neo vgpr_cam ( // @[allocator_neo.scala 129:26]
    .clock(vgpr_cam_clock),
    .reset(vgpr_cam_reset),
    .io_res_search_out(vgpr_cam_io_res_search_out),
    .io_res_search_en(vgpr_cam_io_res_search_en),
    .io_res_search_out_start_0(vgpr_cam_io_res_search_out_start_0),
    .io_res_search_out_start_1(vgpr_cam_io_res_search_out_start_1),
    .io_res_search_size(vgpr_cam_io_res_search_size),
    .io_cam_wr_en(vgpr_cam_io_cam_wr_en),
    .io_cam_wr_addr(vgpr_cam_io_cam_wr_addr),
    .io_cam_wr_data(vgpr_cam_io_cam_wr_data),
    .io_cam_wr_start(vgpr_cam_io_cam_wr_start)
  );
  cam_allocator_neo sgpr_cam ( // @[allocator_neo.scala 130:26]
    .clock(sgpr_cam_clock),
    .reset(sgpr_cam_reset),
    .io_res_search_out(sgpr_cam_io_res_search_out),
    .io_res_search_en(sgpr_cam_io_res_search_en),
    .io_res_search_out_start_0(sgpr_cam_io_res_search_out_start_0),
    .io_res_search_out_start_1(sgpr_cam_io_res_search_out_start_1),
    .io_res_search_size(sgpr_cam_io_res_search_size),
    .io_cam_wr_en(sgpr_cam_io_cam_wr_en),
    .io_cam_wr_addr(sgpr_cam_io_cam_wr_addr),
    .io_cam_wr_data(sgpr_cam_io_cam_wr_data),
    .io_cam_wr_start(sgpr_cam_io_cam_wr_start)
  );
  cam_allocator_neo lds_cam ( // @[allocator_neo.scala 131:25]
    .clock(lds_cam_clock),
    .reset(lds_cam_reset),
    .io_res_search_out(lds_cam_io_res_search_out),
    .io_res_search_en(lds_cam_io_res_search_en),
    .io_res_search_out_start_0(lds_cam_io_res_search_out_start_0),
    .io_res_search_out_start_1(lds_cam_io_res_search_out_start_1),
    .io_res_search_size(lds_cam_io_res_search_size),
    .io_cam_wr_en(lds_cam_io_cam_wr_en),
    .io_cam_wr_addr(lds_cam_io_cam_wr_addr),
    .io_cam_wr_data(lds_cam_io_cam_wr_data),
    .io_cam_wr_start(lds_cam_io_cam_wr_start)
  );
  cam_allocator wf_cam ( // @[allocator_neo.scala 132:24]
    .clock(wf_cam_clock),
    .reset(wf_cam_reset),
    .io_res_search_out(wf_cam_io_res_search_out),
    .io_res_search_en(wf_cam_io_res_search_en),
    .io_res_search_size(wf_cam_io_res_search_size),
    .io_cam_wr_en(wf_cam_io_cam_wr_en),
    .io_cam_wr_addr(wf_cam_io_cam_wr_addr),
    .io_cam_wr_data(wf_cam_io_cam_wr_data)
  );
  cam_allocator wg_cam ( // @[allocator_neo.scala 133:24]
    .clock(wg_cam_clock),
    .reset(wg_cam_reset),
    .io_res_search_out(wg_cam_io_res_search_out),
    .io_res_search_en(wg_cam_io_res_search_en),
    .io_res_search_size(wg_cam_io_res_search_size),
    .io_cam_wr_en(wg_cam_io_cam_wr_en),
    .io_cam_wr_addr(wg_cam_io_cam_wr_addr),
    .io_cam_wr_data(wg_cam_io_cam_wr_data)
  );
  prefer_select prefer_select ( // @[allocator_neo.scala 303:31]
    .io_signal_0(prefer_select_io_signal_0),
    .io_signal_1(prefer_select_io_signal_1),
    .io_prefer(prefer_select_io_prefer),
    .io_valid(prefer_select_io_valid),
    .io_id(prefer_select_io_id)
  );
  assign io_allocator_cu_valid = size_ram_valid; // @[allocator_neo.scala 270:27]
  assign io_allocator_cu_rejected = ~size_ram_cu_id_found; // @[allocator_neo.scala 271:33]
  assign io_allocator_wg_id_out = wg_id_out; // @[allocator_neo.scala 273:28]
  assign io_allocator_cu_id_out = cu_id_out; // @[allocator_neo.scala 272:28]
  assign io_allocator_wf_count = wf_count_out; // @[allocator_neo.scala 274:27]
  assign io_allocator_vgpr_size_out = vgpr_size_out; // @[allocator_neo.scala 276:32]
  assign io_allocator_sgpr_size_out = sgpr_size_out; // @[allocator_neo.scala 277:32]
  assign io_allocator_lds_size_out = lds_size_out; // @[allocator_neo.scala 278:31]
  assign io_allocator_vgpr_start_out = ~_GEN_50 ? 12'h0 : vgpr_start_out; // @[allocator_neo.scala 280:37 281:37 286:37]
  assign io_allocator_sgpr_start_out = ~_GEN_50 ? 12'h0 : sgpr_start_out; // @[allocator_neo.scala 280:37 282:37 287:37]
  assign io_allocator_lds_start_out = ~_GEN_50 ? 12'h0 : lds_start_out; // @[allocator_neo.scala 280:37 283:36 288:36]
  assign vgpr_cam_clock = clock;
  assign vgpr_cam_reset = reset;
  assign vgpr_cam_io_res_search_en = alloc_valid_i; // @[allocator_neo.scala 138:31]
  assign vgpr_cam_io_res_search_size = alloc_vgpr_size_i; // @[allocator_neo.scala 139:33]
  assign vgpr_cam_io_cam_wr_en = cam_up_valid_i; // @[allocator_neo.scala 144:27]
  assign vgpr_cam_io_cam_wr_addr = cam_up_cu_id_i; // @[allocator_neo.scala 145:29]
  assign vgpr_cam_io_cam_wr_data = cam_up_vgpr_size_i; // @[allocator_neo.scala 146:29]
  assign vgpr_cam_io_cam_wr_start = cam_up_vgpr_strt_i; // @[allocator_neo.scala 147:30]
  assign sgpr_cam_clock = clock;
  assign sgpr_cam_reset = reset;
  assign sgpr_cam_io_res_search_en = alloc_valid_i; // @[allocator_neo.scala 149:31]
  assign sgpr_cam_io_res_search_size = alloc_sgpr_size_i; // @[allocator_neo.scala 150:33]
  assign sgpr_cam_io_cam_wr_en = cam_up_valid_i; // @[allocator_neo.scala 155:27]
  assign sgpr_cam_io_cam_wr_addr = cam_up_cu_id_i; // @[allocator_neo.scala 156:29]
  assign sgpr_cam_io_cam_wr_data = cam_up_sgpr_size_i; // @[allocator_neo.scala 157:29]
  assign sgpr_cam_io_cam_wr_start = cam_up_sgpr_strt_i; // @[allocator_neo.scala 158:30]
  assign lds_cam_clock = clock;
  assign lds_cam_reset = reset;
  assign lds_cam_io_res_search_en = alloc_valid_i; // @[allocator_neo.scala 160:30]
  assign lds_cam_io_res_search_size = alloc_lds_size_i; // @[allocator_neo.scala 161:32]
  assign lds_cam_io_cam_wr_en = cam_up_valid_i; // @[allocator_neo.scala 166:26]
  assign lds_cam_io_cam_wr_addr = cam_up_cu_id_i; // @[allocator_neo.scala 167:28]
  assign lds_cam_io_cam_wr_data = cam_up_lds_size_i; // @[allocator_neo.scala 168:28]
  assign lds_cam_io_cam_wr_start = cam_up_lds_strt_i; // @[allocator_neo.scala 169:29]
  assign wf_cam_clock = clock;
  assign wf_cam_reset = reset;
  assign wf_cam_io_res_search_en = alloc_valid_i; // @[allocator_neo.scala 171:29]
  assign wf_cam_io_res_search_size = {{1'd0}, alloc_num_wf_i}; // @[allocator_neo.scala 173:31]
  assign wf_cam_io_cam_wr_en = cam_up_valid_i; // @[allocator_neo.scala 177:25]
  assign wf_cam_io_cam_wr_addr = cam_up_cu_id_i; // @[allocator_neo.scala 178:27]
  assign wf_cam_io_cam_wr_data = {{1'd0}, cam_up_wf_count_i}; // @[allocator_neo.scala 179:27]
  assign wg_cam_clock = clock;
  assign wg_cam_reset = reset;
  assign wg_cam_io_res_search_en = alloc_valid_i; // @[allocator_neo.scala 181:29]
  assign wg_cam_io_res_search_size = 4'h1; // @[allocator_neo.scala 182:31]
  assign wg_cam_io_cam_wr_en = cam_up_valid_i; // @[allocator_neo.scala 184:25]
  assign wg_cam_io_cam_wr_addr = cam_up_cu_id_i; // @[allocator_neo.scala 185:27]
  assign wg_cam_io_cam_wr_data = {{1'd0}, cam_up_wg_count_i}; // @[allocator_neo.scala 186:27]
  assign prefer_select_io_signal_0 = anded_cam_out[0]; // @[allocator_neo.scala 304:46]
  assign prefer_select_io_signal_1 = anded_cam_out[1]; // @[allocator_neo.scala 304:46]
  assign prefer_select_io_prefer = anded_cam_wg_id[1:0]; // @[allocator_neo.scala 305:47]
  always @(posedge clock) begin
    if (reset) begin // @[allocator_neo.scala 42:32]
      alloc_valid_i <= 1'h0; // @[allocator_neo.scala 42:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      alloc_valid_i <= io_dis_controller_start_alloc; // @[allocator_neo.scala 202:23]
    end
    if (reset) begin // @[allocator_neo.scala 43:32]
      alloc_wg_id_i <= 5'h0; // @[allocator_neo.scala 43:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      alloc_wg_id_i <= io_inflight_wg_buffer_alloc_wg_id; // @[allocator_neo.scala 203:23]
    end
    if (reset) begin // @[allocator_neo.scala 44:33]
      alloc_num_wf_i <= 3'h0; // @[allocator_neo.scala 44:33]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      alloc_num_wf_i <= io_inflight_wg_buffer_alloc_num_wf; // @[allocator_neo.scala 204:24]
    end
    if (reset) begin // @[allocator_neo.scala 45:36]
      alloc_vgpr_size_i <= 13'h0; // @[allocator_neo.scala 45:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      alloc_vgpr_size_i <= io_inflight_wg_buffer_alloc_vgpr_size; // @[allocator_neo.scala 205:27]
    end
    if (reset) begin // @[allocator_neo.scala 46:36]
      alloc_sgpr_size_i <= 13'h0; // @[allocator_neo.scala 46:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      alloc_sgpr_size_i <= io_inflight_wg_buffer_alloc_sgpr_size; // @[allocator_neo.scala 206:27]
    end
    if (reset) begin // @[allocator_neo.scala 47:35]
      alloc_lds_size_i <= 13'h0; // @[allocator_neo.scala 47:35]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      alloc_lds_size_i <= io_inflight_wg_buffer_alloc_lds_size; // @[allocator_neo.scala 207:26]
    end
    if (reset) begin // @[allocator_neo.scala 48:43]
      dis_controller_cu_busy_i <= 2'h0; // @[allocator_neo.scala 48:43]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      dis_controller_cu_busy_i <= io_dis_controller_cu_busy; // @[allocator_neo.scala 208:34]
    end
    if (reset) begin // @[allocator_neo.scala 50:33]
      cam_up_valid_i <= 1'h0; // @[allocator_neo.scala 50:33]
    end else begin
      cam_up_valid_i <= io_grt_cam_up_valid; // @[allocator_neo.scala 256:20]
    end
    if (reset) begin // @[allocator_neo.scala 51:33]
      cam_up_cu_id_i <= 2'h0; // @[allocator_neo.scala 51:33]
    end else begin
      cam_up_cu_id_i <= io_grt_cam_up_cu_id; // @[allocator_neo.scala 257:20]
    end
    if (reset) begin // @[allocator_neo.scala 52:37]
      cam_up_vgpr_strt_i <= 12'h0; // @[allocator_neo.scala 52:37]
    end else begin
      cam_up_vgpr_strt_i <= io_grt_cam_up_vgpr_strt; // @[allocator_neo.scala 260:24]
    end
    if (reset) begin // @[allocator_neo.scala 53:37]
      cam_up_vgpr_size_i <= 13'h0; // @[allocator_neo.scala 53:37]
    end else begin
      cam_up_vgpr_size_i <= io_grt_cam_up_vgpr_size; // @[allocator_neo.scala 267:24]
    end
    if (reset) begin // @[allocator_neo.scala 54:37]
      cam_up_sgpr_strt_i <= 12'h0; // @[allocator_neo.scala 54:37]
    end else begin
      cam_up_sgpr_strt_i <= io_grt_cam_up_sgpr_strt; // @[allocator_neo.scala 261:24]
    end
    if (reset) begin // @[allocator_neo.scala 55:37]
      cam_up_sgpr_size_i <= 13'h0; // @[allocator_neo.scala 55:37]
    end else begin
      cam_up_sgpr_size_i <= io_grt_cam_up_sgpr_size; // @[allocator_neo.scala 268:24]
    end
    if (reset) begin // @[allocator_neo.scala 56:36]
      cam_up_lds_strt_i <= 12'h0; // @[allocator_neo.scala 56:36]
    end else begin
      cam_up_lds_strt_i <= io_grt_cam_up_lds_strt; // @[allocator_neo.scala 262:23]
    end
    if (reset) begin // @[allocator_neo.scala 57:36]
      cam_up_lds_size_i <= 13'h0; // @[allocator_neo.scala 57:36]
    end else begin
      cam_up_lds_size_i <= io_grt_cam_up_lds_size; // @[allocator_neo.scala 266:23]
    end
    if (reset) begin // @[allocator_neo.scala 58:36]
      cam_up_wf_count_i <= 3'h0; // @[allocator_neo.scala 58:36]
    end else begin
      cam_up_wf_count_i <= io_grt_cam_up_wf_count; // @[allocator_neo.scala 258:23]
    end
    if (reset) begin // @[allocator_neo.scala 59:36]
      cam_up_wg_count_i <= 3'h0; // @[allocator_neo.scala 59:36]
    end else begin
      cam_up_wg_count_i <= io_grt_cam_up_wg_count; // @[allocator_neo.scala 259:23]
    end
    if (reset) begin // @[allocator_neo.scala 70:33]
      cam_wait_valid <= 1'h0; // @[allocator_neo.scala 70:33]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_valid <= alloc_valid_i; // @[allocator_neo.scala 211:24]
    end
    if (reset) begin // @[allocator_neo.scala 71:33]
      cam_wait_wg_id <= 5'h0; // @[allocator_neo.scala 71:33]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_wg_id <= alloc_wg_id_i; // @[allocator_neo.scala 212:24]
    end
    if (reset) begin // @[allocator_neo.scala 72:36]
      cam_wait_wf_count <= 3'h0; // @[allocator_neo.scala 72:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_wf_count <= alloc_num_wf_i; // @[allocator_neo.scala 213:27]
    end
    if (reset) begin // @[allocator_neo.scala 73:37]
      cam_wait_vgpr_size <= 13'h0; // @[allocator_neo.scala 73:37]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_vgpr_size <= alloc_vgpr_size_i; // @[allocator_neo.scala 214:28]
    end
    if (reset) begin // @[allocator_neo.scala 74:37]
      cam_wait_sgpr_size <= 13'h0; // @[allocator_neo.scala 74:37]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_sgpr_size <= alloc_sgpr_size_i; // @[allocator_neo.scala 215:28]
    end
    if (reset) begin // @[allocator_neo.scala 75:36]
      cam_wait_lds_size <= 13'h0; // @[allocator_neo.scala 75:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_lds_size <= alloc_lds_size_i; // @[allocator_neo.scala 216:27]
    end
    if (reset) begin // @[allocator_neo.scala 76:50]
      cam_wait_dis_controller_cu_busy <= 2'h0; // @[allocator_neo.scala 76:50]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cam_wait_dis_controller_cu_busy <= dis_controller_cu_busy_i; // @[allocator_neo.scala 217:41]
    end
    if (reset) begin // @[allocator_neo.scala 79:38]
      anded_cam_out_valid <= 1'h0; // @[allocator_neo.scala 79:38]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_out_valid <= cam_wait_valid; // @[allocator_neo.scala 220:29]
    end
    if (reset) begin // @[allocator_neo.scala 80:32]
      anded_cam_out <= 2'h0; // @[allocator_neo.scala 80:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_out <= _anded_cam_out_T_5; // @[allocator_neo.scala 221:23]
    end
    if (reset) begin // @[allocator_neo.scala 81:34]
      anded_cam_wg_id <= 5'h0; // @[allocator_neo.scala 81:34]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_wg_id <= cam_wait_wg_id; // @[allocator_neo.scala 222:25]
    end
    if (reset) begin // @[allocator_neo.scala 82:37]
      anded_cam_wf_count <= 3'h0; // @[allocator_neo.scala 82:37]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_wf_count <= cam_wait_wf_count; // @[allocator_neo.scala 223:28]
    end
    if (reset) begin // @[allocator_neo.scala 83:38]
      anded_cam_vgpr_size <= 13'h0; // @[allocator_neo.scala 83:38]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_vgpr_size <= cam_wait_vgpr_size; // @[allocator_neo.scala 224:29]
    end
    if (reset) begin // @[allocator_neo.scala 84:38]
      anded_cam_sgpr_size <= 13'h0; // @[allocator_neo.scala 84:38]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_sgpr_size <= cam_wait_sgpr_size; // @[allocator_neo.scala 225:29]
    end
    if (reset) begin // @[allocator_neo.scala 85:37]
      anded_cam_lds_size <= 13'h0; // @[allocator_neo.scala 85:37]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      anded_cam_lds_size <= cam_wait_lds_size; // @[allocator_neo.scala 226:28]
    end
    if (reset) begin // @[allocator_neo.scala 88:39]
      encoded_cu_out_valid <= 1'h0; // @[allocator_neo.scala 88:39]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_cu_out_valid <= anded_cam_out_valid; // @[allocator_neo.scala 229:30]
    end
    if (reset) begin // @[allocator_neo.scala 89:41]
      encoded_cu_found_valid <= 1'h0; // @[allocator_neo.scala 89:41]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_cu_found_valid <= encoded_cu_found_valid_comb; // @[allocator_neo.scala 230:32]
    end
    if (reset) begin // @[allocator_neo.scala 91:32]
      encoded_cu_id <= 2'h0; // @[allocator_neo.scala 91:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_cu_id <= encoded_cu_id_comb; // @[allocator_neo.scala 231:23]
    end
    if (reset) begin // @[allocator_neo.scala 93:35]
      encoded_cu_wg_id <= 5'h0; // @[allocator_neo.scala 93:35]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_cu_wg_id <= anded_cam_wg_id; // @[allocator_neo.scala 233:26]
    end
    if (reset) begin // @[allocator_neo.scala 94:35]
      encoded_wf_count <= 3'h0; // @[allocator_neo.scala 94:35]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_wf_count <= anded_cam_wf_count; // @[allocator_neo.scala 232:26]
    end
    if (reset) begin // @[allocator_neo.scala 95:36]
      encoded_vgpr_size <= 13'h0; // @[allocator_neo.scala 95:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_vgpr_size <= anded_cam_vgpr_size; // @[allocator_neo.scala 234:27]
    end
    if (reset) begin // @[allocator_neo.scala 96:36]
      encoded_sgpr_size <= 13'h0; // @[allocator_neo.scala 96:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_sgpr_size <= anded_cam_sgpr_size; // @[allocator_neo.scala 235:27]
    end
    if (reset) begin // @[allocator_neo.scala 97:35]
      encoded_lds_size <= 13'h0; // @[allocator_neo.scala 97:35]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      encoded_lds_size <= anded_cam_lds_size; // @[allocator_neo.scala 236:26]
    end
    if (reset) begin // @[allocator_neo.scala 98:37]
      encoded_vgpr_start <= 12'h0; // @[allocator_neo.scala 98:37]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      if (encoded_cu_id_comb[0]) begin // @[allocator_neo.scala 308:29]
        encoded_vgpr_start <= vgpr_cam_start_vec_1; // @[allocator_neo.scala 308:29]
      end else begin
        encoded_vgpr_start <= vgpr_cam_start_vec_0;
      end
    end
    if (reset) begin // @[allocator_neo.scala 99:37]
      encoded_sgpr_start <= 12'h0; // @[allocator_neo.scala 99:37]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      if (encoded_cu_id_comb[0]) begin // @[allocator_neo.scala 307:29]
        encoded_sgpr_start <= sgpr_cam_start_vec_1; // @[allocator_neo.scala 307:29]
      end else begin
        encoded_sgpr_start <= sgpr_cam_start_vec_0;
      end
    end
    if (reset) begin // @[allocator_neo.scala 100:36]
      encoded_lds_start <= 12'h0; // @[allocator_neo.scala 100:36]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      if (encoded_cu_id_comb[0]) begin // @[allocator_neo.scala 309:28]
        encoded_lds_start <= lds_cam_start_vec_1; // @[allocator_neo.scala 309:28]
      end else begin
        encoded_lds_start <= lds_cam_start_vec_0;
      end
    end
    if (reset) begin // @[allocator_neo.scala 103:33]
      size_ram_valid <= 1'h0; // @[allocator_neo.scala 103:33]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      size_ram_valid <= encoded_cu_out_valid; // @[allocator_neo.scala 243:24]
    end
    if (reset) begin // @[allocator_neo.scala 104:39]
      size_ram_cu_id_found <= 1'h0; // @[allocator_neo.scala 104:39]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      size_ram_cu_id_found <= encoded_cu_found_valid; // @[allocator_neo.scala 244:30]
    end
    if (reset) begin // @[allocator_neo.scala 105:28]
      cu_id_out <= 2'h0; // @[allocator_neo.scala 105:28]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      cu_id_out <= encoded_cu_id; // @[allocator_neo.scala 245:19]
    end
    if (reset) begin // @[allocator_neo.scala 106:33]
      vgpr_start_out <= 12'h0; // @[allocator_neo.scala 106:33]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      vgpr_start_out <= encoded_vgpr_start; // @[allocator_neo.scala 252:24]
    end
    if (reset) begin // @[allocator_neo.scala 107:33]
      sgpr_start_out <= 12'h0; // @[allocator_neo.scala 107:33]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      sgpr_start_out <= encoded_sgpr_start; // @[allocator_neo.scala 253:24]
    end
    if (reset) begin // @[allocator_neo.scala 108:32]
      lds_start_out <= 12'h0; // @[allocator_neo.scala 108:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      lds_start_out <= encoded_lds_start; // @[allocator_neo.scala 251:23]
    end
    if (reset) begin // @[allocator_neo.scala 109:28]
      wg_id_out <= 5'h0; // @[allocator_neo.scala 109:28]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      wg_id_out <= encoded_cu_wg_id; // @[allocator_neo.scala 247:19]
    end
    if (reset) begin // @[allocator_neo.scala 110:31]
      wf_count_out <= 3'h0; // @[allocator_neo.scala 110:31]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      wf_count_out <= encoded_wf_count; // @[allocator_neo.scala 246:22]
    end
    if (reset) begin // @[allocator_neo.scala 111:32]
      vgpr_size_out <= 13'h0; // @[allocator_neo.scala 111:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      vgpr_size_out <= encoded_vgpr_size; // @[allocator_neo.scala 248:23]
    end
    if (reset) begin // @[allocator_neo.scala 112:32]
      sgpr_size_out <= 13'h0; // @[allocator_neo.scala 112:32]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      sgpr_size_out <= encoded_sgpr_size; // @[allocator_neo.scala 249:23]
    end
    if (reset) begin // @[allocator_neo.scala 113:31]
      lds_size_out <= 13'h0; // @[allocator_neo.scala 113:31]
    end else if (_T) begin // @[allocator_neo.scala 200:28]
      lds_size_out <= encoded_lds_size; // @[allocator_neo.scala 250:22]
    end
    if (reset) begin // @[allocator_neo.scala 125:33]
      cu_initialized_0 <= 1'h0; // @[allocator_neo.scala 125:33]
    end else if (cam_up_valid_i) begin // @[allocator_neo.scala 263:25]
      cu_initialized_0 <= _GEN_45;
    end
    if (reset) begin // @[allocator_neo.scala 125:33]
      cu_initialized_1 <= 1'h0; // @[allocator_neo.scala 125:33]
    end else if (cam_up_valid_i) begin // @[allocator_neo.scala 263:25]
      cu_initialized_1 <= _GEN_46;
    end
    if (reset) begin // @[allocator_neo.scala 127:35]
      pipeline_waiting <= 1'h0; // @[allocator_neo.scala 127:35]
    end else if (io_dis_controller_alloc_ack) begin // @[allocator_neo.scala 196:38]
      pipeline_waiting <= 1'h0; // @[allocator_neo.scala 197:26]
    end else begin
      pipeline_waiting <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  alloc_valid_i = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  alloc_wg_id_i = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  alloc_num_wf_i = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  alloc_vgpr_size_i = _RAND_3[12:0];
  _RAND_4 = {1{`RANDOM}};
  alloc_sgpr_size_i = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  alloc_lds_size_i = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  dis_controller_cu_busy_i = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  cam_up_valid_i = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cam_up_cu_id_i = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  cam_up_vgpr_strt_i = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  cam_up_vgpr_size_i = _RAND_10[12:0];
  _RAND_11 = {1{`RANDOM}};
  cam_up_sgpr_strt_i = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  cam_up_sgpr_size_i = _RAND_12[12:0];
  _RAND_13 = {1{`RANDOM}};
  cam_up_lds_strt_i = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  cam_up_lds_size_i = _RAND_14[12:0];
  _RAND_15 = {1{`RANDOM}};
  cam_up_wf_count_i = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  cam_up_wg_count_i = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  cam_wait_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  cam_wait_wg_id = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  cam_wait_wf_count = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  cam_wait_vgpr_size = _RAND_20[12:0];
  _RAND_21 = {1{`RANDOM}};
  cam_wait_sgpr_size = _RAND_21[12:0];
  _RAND_22 = {1{`RANDOM}};
  cam_wait_lds_size = _RAND_22[12:0];
  _RAND_23 = {1{`RANDOM}};
  cam_wait_dis_controller_cu_busy = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  anded_cam_out_valid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  anded_cam_out = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  anded_cam_wg_id = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  anded_cam_wf_count = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  anded_cam_vgpr_size = _RAND_28[12:0];
  _RAND_29 = {1{`RANDOM}};
  anded_cam_sgpr_size = _RAND_29[12:0];
  _RAND_30 = {1{`RANDOM}};
  anded_cam_lds_size = _RAND_30[12:0];
  _RAND_31 = {1{`RANDOM}};
  encoded_cu_out_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  encoded_cu_found_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  encoded_cu_id = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  encoded_cu_wg_id = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  encoded_wf_count = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  encoded_vgpr_size = _RAND_36[12:0];
  _RAND_37 = {1{`RANDOM}};
  encoded_sgpr_size = _RAND_37[12:0];
  _RAND_38 = {1{`RANDOM}};
  encoded_lds_size = _RAND_38[12:0];
  _RAND_39 = {1{`RANDOM}};
  encoded_vgpr_start = _RAND_39[11:0];
  _RAND_40 = {1{`RANDOM}};
  encoded_sgpr_start = _RAND_40[11:0];
  _RAND_41 = {1{`RANDOM}};
  encoded_lds_start = _RAND_41[11:0];
  _RAND_42 = {1{`RANDOM}};
  size_ram_valid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  size_ram_cu_id_found = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  cu_id_out = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  vgpr_start_out = _RAND_45[11:0];
  _RAND_46 = {1{`RANDOM}};
  sgpr_start_out = _RAND_46[11:0];
  _RAND_47 = {1{`RANDOM}};
  lds_start_out = _RAND_47[11:0];
  _RAND_48 = {1{`RANDOM}};
  wg_id_out = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  wf_count_out = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  vgpr_size_out = _RAND_50[12:0];
  _RAND_51 = {1{`RANDOM}};
  sgpr_size_out = _RAND_51[12:0];
  _RAND_52 = {1{`RANDOM}};
  lds_size_out = _RAND_52[12:0];
  _RAND_53 = {1{`RANDOM}};
  cu_initialized_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  cu_initialized_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  pipeline_waiting = _RAND_55[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module resource_table(
  input         clock,
  input         reset,
  output        io_res_table_done_o,
  output [13:0] io_cam_biggest_space_size,
  output [12:0] io_cam_biggest_space_addr,
  input         io_alloc_res_en,
  input         io_dealloc_res_en,
  input         io_alloc_cu_id,
  input         io_dealloc_cu_id,
  input  [1:0]  io_alloc_wg_slot_id,
  input  [1:0]  io_dealloc_wg_slot_id,
  input  [13:0] io_alloc_res_size,
  input  [12:0] io_alloc_res_start
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
`endif // RANDOMIZE_REG_INIT
  reg  res_table_done; // @[resource_table.scala 24:33]
  reg  alloc_res_en_i; // @[resource_table.scala 39:33]
  reg  dealloc_res_en_i; // @[resource_table.scala 40:35]
  reg [1:0] alloc_wg_slot_id_i; // @[resource_table.scala 43:37]
  reg [1:0] dealloc_wg_slot_id_i; // @[resource_table.scala 44:39]
  reg [13:0] alloc_res_size_i; // @[resource_table.scala 46:35]
  reg [12:0] alloc_res_start_i; // @[resource_table.scala 47:36]
  reg [30:0] resource_table_ram_0; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_1; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_2; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_3; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_4; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_5; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_6; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_7; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_8; // @[resource_table.scala 80:37]
  reg [30:0] resource_table_ram_9; // @[resource_table.scala 80:37]
  reg [1:0] table_head_pointer_0; // @[resource_table.scala 81:37]
  reg [1:0] table_head_pointer_1; // @[resource_table.scala 81:37]
  reg [1:0] table_head_pointer_i; // @[resource_table.scala 82:39]
  reg [3:0] m_state; // @[resource_table.scala 103:26]
  reg [3:0] a_state; // @[resource_table.scala 110:26]
  reg [4:0] d_state; // @[resource_table.scala 118:26]
  reg [3:0] f_state; // @[resource_table.scala 126:26]
  reg [30:0] res_table_wr_reg; // @[resource_table.scala 129:35]
  reg [30:0] res_table_rd_reg; // @[resource_table.scala 130:35]
  reg [30:0] res_table_last_rd_reg; // @[resource_table.scala 131:40]
  reg  res_addr_cu_id; // @[resource_table.scala 132:33]
  reg [1:0] res_addr_wg_slot; // @[resource_table.scala 133:35]
  reg  res_table_rd_en; // @[resource_table.scala 134:34]
  reg  res_table_wr_en; // @[resource_table.scala 135:34]
  reg  res_table_rd_valid; // @[resource_table.scala 136:37]
  reg [13:0] res_table_max_size; // @[resource_table.scala 137:37]
  reg [12:0] res_table_max_start; // @[resource_table.scala 138:38]
  reg  alloc_start; // @[resource_table.scala 141:30]
  reg  dealloc_start; // @[resource_table.scala 142:32]
  reg  find_max_start; // @[resource_table.scala 143:33]
  reg  alloc_done; // @[resource_table.scala 144:29]
  reg  dealloc_done; // @[resource_table.scala 145:31]
  reg  find_max_done; // @[resource_table.scala 146:32]
  reg  new_entry_is_last; // @[resource_table.scala 147:36]
  reg  new_entry_is_first; // @[resource_table.scala 148:37]
  reg  rem_entry_is_last; // @[resource_table.scala 149:36]
  reg  rem_entry_is_first; // @[resource_table.scala 150:37]
  reg  cu_initialized_0; // @[resource_table.scala 151:33]
  reg  cu_initialized_1; // @[resource_table.scala 151:33]
  reg  cu_initialized_i; // @[resource_table.scala 152:35]
  wire [12:0] rtrr_res_strt = res_table_rd_reg[12:0]; // @[resource_table.scala 59:20]
  wire [12:0] rtlrr_res_strt = res_table_last_rd_reg[12:0]; // @[resource_table.scala 59:20]
  wire [13:0] rtrr_res_size = res_table_rd_reg[26:13]; // @[resource_table.scala 62:20]
  wire [13:0] rtlrr_res_size = res_table_last_rd_reg[26:13]; // @[resource_table.scala 62:20]
  wire  _GEN_12 = alloc_res_en_i ? 1'h0 : dealloc_res_en_i; // @[resource_table.scala 187:19 192:33]
  wire [3:0] _GEN_16 = dealloc_done ? 4'h8 : m_state; // @[resource_table.scala 208:31 210:25 103:26]
  wire [3:0] _GEN_18 = find_max_done ? 4'h1 : m_state; // @[resource_table.scala 214:32 216:25 103:26]
  wire [3:0] _GEN_20 = 4'h8 == m_state ? _GEN_18 : m_state; // @[resource_table.scala 190:20 103:26]
  wire  _GEN_21 = 4'h4 == m_state & dealloc_done; // @[resource_table.scala 188:20 190:20]
  wire  _GEN_27 = 4'h1 == m_state & alloc_res_en_i; // @[resource_table.scala 186:17 190:20]
  wire  _GEN_29 = 4'h1 == m_state & _GEN_12; // @[resource_table.scala 187:19 190:20]
  wire  _T_5 = table_head_pointer_i == 2'h3; // @[resource_table.scala 235:43]
  wire  _T_7 = table_head_pointer_i == 2'h3 | ~cu_initialized_i; // @[resource_table.scala 235:69]
  wire  _GEN_34 = table_head_pointer_i == 2'h3 | ~cu_initialized_i ? 1'h0 : 1'h1; // @[resource_table.scala 224:21 235:90 243:37]
  wire [1:0] _GEN_35 = table_head_pointer_i == 2'h3 | ~cu_initialized_i ? res_addr_wg_slot : table_head_pointer_i; // @[resource_table.scala 133:35 235:90 244:38]
  wire  _GEN_39 = alloc_start & _GEN_34; // @[resource_table.scala 224:21 230:30]
  wire [1:0] _GEN_40 = alloc_start ? _GEN_35 : res_addr_wg_slot; // @[resource_table.scala 230:30 133:35]
  wire  _T_12 = res_table_rd_reg[28:27] == 2'h2; // @[resource_table.scala 255:66]
  wire [30:0] _res_table_wr_reg_T_3 = {res_table_rd_reg[30:29],alloc_wg_slot_id_i,rtrr_res_size,rtrr_res_strt}; // @[Cat.scala 31:58]
  wire  _GEN_41 = res_table_rd_reg[28:27] == 2'h2 | new_entry_is_first; // @[resource_table.scala 148:37 255:95 256:44]
  wire [30:0] _GEN_43 = res_table_rd_reg[28:27] == 2'h2 ? _res_table_wr_reg_T_3 : _res_table_wr_reg_T_3; // @[resource_table.scala 255:95 258:42 263:42]
  wire [3:0] _GEN_44 = res_table_rd_reg[28:27] == 2'h2 ? 4'h8 : 4'h4; // @[resource_table.scala 255:95 259:33 264:33]
  wire  _T_14 = res_table_rd_reg[30:29] == 2'h3; // @[resource_table.scala 267:67]
  wire [30:0] _res_table_wr_reg_T_11 = {alloc_wg_slot_id_i,res_table_rd_reg[28:27],rtrr_res_size,rtrr_res_strt}; // @[Cat.scala 31:58]
  wire [30:0] _GEN_46 = res_table_rd_reg[30:29] == 2'h3 ? _res_table_wr_reg_T_11 : res_table_wr_reg; // @[resource_table.scala 129:35 267:93 270:38]
  wire  _GEN_47 = res_table_rd_reg[30:29] == 2'h3 | new_entry_is_last; // @[resource_table.scala 147:36 267:93 271:39]
  wire [3:0] _GEN_48 = res_table_rd_reg[30:29] == 2'h3 ? 4'h8 : a_state; // @[resource_table.scala 110:26 267:93 272:29]
  wire  _GEN_49 = res_table_rd_reg[30:29] == 2'h3 ? 1'h0 : 1'h1; // @[resource_table.scala 224:21 267:93 276:37]
  wire [1:0] _GEN_50 = res_table_rd_reg[30:29] == 2'h3 ? res_addr_wg_slot : res_table_rd_reg[30:29]; // @[resource_table.scala 133:35 267:93 277:38]
  wire  _GEN_51 = rtrr_res_strt > alloc_res_start_i ? _GEN_41 : new_entry_is_first; // @[resource_table.scala 148:37 253:74]
  wire  _GEN_52 = rtrr_res_strt > alloc_res_start_i | _T_14; // @[resource_table.scala 253:74]
  wire [30:0] _GEN_53 = rtrr_res_strt > alloc_res_start_i ? _GEN_43 : _GEN_46; // @[resource_table.scala 253:74]
  wire [3:0] _GEN_54 = rtrr_res_strt > alloc_res_start_i ? _GEN_44 : _GEN_48; // @[resource_table.scala 253:74]
  wire  _GEN_55 = rtrr_res_strt > alloc_res_start_i ? new_entry_is_last : _GEN_47; // @[resource_table.scala 147:36 253:74]
  wire  _GEN_56 = rtrr_res_strt > alloc_res_start_i ? 1'h0 : _GEN_49; // @[resource_table.scala 224:21 253:74]
  wire [1:0] _GEN_57 = rtrr_res_strt > alloc_res_start_i ? res_addr_wg_slot : _GEN_50; // @[resource_table.scala 133:35 253:74]
  wire  _GEN_59 = res_table_rd_valid & _GEN_52; // @[resource_table.scala 225:21 251:37]
  wire [30:0] _GEN_60 = res_table_rd_valid ? _GEN_53 : res_table_wr_reg; // @[resource_table.scala 129:35 251:37]
  wire  _GEN_63 = res_table_rd_valid & _GEN_56; // @[resource_table.scala 224:21 251:37]
  wire [1:0] _GEN_64 = res_table_rd_valid ? _GEN_57 : res_addr_wg_slot; // @[resource_table.scala 133:35 251:37]
  wire [30:0] _res_table_wr_reg_T_15 = {alloc_wg_slot_id_i,res_table_last_rd_reg[28:27],rtlrr_res_size,rtlrr_res_strt}; // @[Cat.scala 31:58]
  wire [1:0] _GEN_65 = new_entry_is_first ? alloc_wg_slot_id_i : table_head_pointer_i; // @[resource_table.scala 289:37 290:38 82:39]
  wire [30:0] _res_table_wr_reg_T_16 = {4'he,alloc_res_size_i,alloc_res_start_i}; // @[Cat.scala 31:58]
  wire [30:0] _res_table_wr_reg_T_17 = {2'h3,res_addr_wg_slot,alloc_res_size_i,alloc_res_start_i}; // @[Cat.scala 31:58]
  wire [30:0] _res_table_wr_reg_T_18 = {res_addr_wg_slot,2'h2,alloc_res_size_i,alloc_res_start_i}; // @[Cat.scala 31:58]
  wire [30:0] _res_table_wr_reg_T_20 = {res_table_last_rd_reg[30:29],res_addr_wg_slot,alloc_res_size_i,alloc_res_start_i
    }; // @[Cat.scala 31:58]
  wire [30:0] _GEN_66 = new_entry_is_first ? _res_table_wr_reg_T_18 : _res_table_wr_reg_T_20; // @[resource_table.scala 303:42 304:34 307:34]
  wire [30:0] _GEN_67 = new_entry_is_last ? _res_table_wr_reg_T_17 : _GEN_66; // @[resource_table.scala 300:41 301:34]
  wire [30:0] _GEN_68 = new_entry_is_first & new_entry_is_last ? _res_table_wr_reg_T_16 : _GEN_67; // @[resource_table.scala 297:58 298:34]
  wire [1:0] _GEN_69 = 4'h8 == a_state ? _GEN_65 : table_head_pointer_i; // @[resource_table.scala 228:20 82:39]
  wire [1:0] _GEN_71 = 4'h8 == a_state ? alloc_wg_slot_id_i : res_addr_wg_slot; // @[resource_table.scala 228:20 295:30 133:35]
  wire [30:0] _GEN_72 = 4'h8 == a_state ? _GEN_68 : res_table_wr_reg; // @[resource_table.scala 228:20 129:35]
  wire [3:0] _GEN_73 = 4'h8 == a_state ? 4'h1 : a_state; // @[resource_table.scala 228:20 310:21 110:26]
  wire  _GEN_74 = 4'h4 == a_state | 4'h8 == a_state; // @[resource_table.scala 228:20 283:29]
  wire [30:0] _GEN_75 = 4'h4 == a_state ? _res_table_wr_reg_T_15 : _GEN_72; // @[resource_table.scala 228:20 284:30]
  wire [1:0] _GEN_76 = 4'h4 == a_state ? res_table_rd_reg[28:27] : _GEN_71; // @[resource_table.scala 228:20 285:30]
  wire [1:0] _GEN_78 = 4'h4 == a_state ? table_head_pointer_i : _GEN_69; // @[resource_table.scala 228:20 82:39]
  wire  _GEN_81 = 4'h2 == a_state ? _GEN_59 : _GEN_74; // @[resource_table.scala 228:20]
  wire [30:0] _GEN_82 = 4'h2 == a_state ? _GEN_60 : _GEN_75; // @[resource_table.scala 228:20]
  wire  _GEN_85 = 4'h2 == a_state & _GEN_63; // @[resource_table.scala 228:20 224:21]
  wire [1:0] _GEN_86 = 4'h2 == a_state ? _GEN_64 : _GEN_76; // @[resource_table.scala 228:20]
  wire [1:0] _GEN_87 = 4'h2 == a_state ? table_head_pointer_i : _GEN_78; // @[resource_table.scala 228:20 82:39]
  wire  _GEN_92 = 4'h1 == a_state ? _GEN_39 : _GEN_85; // @[resource_table.scala 228:20]
  wire [1:0] _GEN_93 = 4'h1 == a_state ? _GEN_40 : _GEN_86; // @[resource_table.scala 228:20]
  wire  _GEN_94 = 4'h1 == a_state ? 1'h0 : _GEN_81; // @[resource_table.scala 228:20 225:21]
  wire [30:0] _GEN_95 = 4'h1 == a_state ? res_table_wr_reg : _GEN_82; // @[resource_table.scala 228:20 129:35]
  wire [1:0] _GEN_96 = 4'h1 == a_state ? table_head_pointer_i : _GEN_87; // @[resource_table.scala 228:20 82:39]
  wire  _GEN_100 = dealloc_start | _GEN_92; // @[resource_table.scala 317:32 320:33]
  wire [1:0] _GEN_101 = dealloc_start ? dealloc_wg_slot_id_i : _GEN_93; // @[resource_table.scala 317:32 321:34]
  wire  _T_24 = _T_12 & _T_14; // @[resource_table.scala 329:91]
  wire  _GEN_103 = _T_14 | rem_entry_is_last; // @[resource_table.scala 149:36 340:93 341:39]
  wire [1:0] _GEN_105 = _T_14 ? res_table_rd_reg[28:27] : res_table_rd_reg[28:27]; // @[resource_table.scala 340:93 343:38 349:38]
  wire [3:0] _GEN_106 = _T_14 ? 4'h8 : 4'h4; // @[resource_table.scala 340:93 344:29 350:29]
  wire  _GEN_107 = _T_12 | rem_entry_is_first; // @[resource_table.scala 150:37 335:96 336:40]
  wire [3:0] _GEN_108 = _T_12 ? 4'h4 : _GEN_106; // @[resource_table.scala 335:96 337:29]
  wire  _GEN_109 = _T_12 ? rem_entry_is_last : _GEN_103; // @[resource_table.scala 149:36 335:96]
  wire  _GEN_110 = _T_12 ? _GEN_92 : 1'h1; // @[resource_table.scala 335:96]
  wire [1:0] _GEN_111 = _T_12 ? _GEN_93 : _GEN_105; // @[resource_table.scala 335:96]
  wire [1:0] _GEN_112 = _T_12 & _T_14 ? 2'h3 : _GEN_96; // @[resource_table.scala 329:160 330:42]
  wire [3:0] _GEN_114 = _T_12 & _T_14 ? 4'h1 : _GEN_108; // @[resource_table.scala 329:160 332:29]
  wire  _GEN_115 = _T_12 & _T_14 ? rem_entry_is_first : _GEN_107; // @[resource_table.scala 329:160 150:37]
  wire  _GEN_116 = _T_12 & _T_14 ? rem_entry_is_last : _GEN_109; // @[resource_table.scala 329:160 149:36]
  wire  _GEN_117 = _T_12 & _T_14 ? _GEN_92 : _GEN_110; // @[resource_table.scala 329:160]
  wire [1:0] _GEN_118 = _T_12 & _T_14 ? _GEN_93 : _GEN_111; // @[resource_table.scala 329:160]
  wire [1:0] _GEN_119 = res_table_rd_valid ? _GEN_112 : _GEN_96; // @[resource_table.scala 327:37]
  wire  _GEN_120 = res_table_rd_valid & _T_24; // @[resource_table.scala 314:18 327:37]
  wire  _GEN_124 = res_table_rd_valid ? _GEN_117 : _GEN_92; // @[resource_table.scala 327:37]
  wire [1:0] _GEN_125 = res_table_rd_valid ? _GEN_118 : _GEN_93; // @[resource_table.scala 327:37]
  wire [30:0] _res_table_wr_reg_T_24 = {res_addr_wg_slot,res_table_rd_reg[28:27],rtrr_res_size,rtrr_res_strt}; // @[Cat.scala 31:58]
  wire [1:0] _GEN_127 = rem_entry_is_last ? _GEN_93 : res_table_last_rd_reg[28:27]; // @[resource_table.scala 367:41 371:34]
  wire  _GEN_128 = rem_entry_is_last ? _GEN_94 : 1'h1; // @[resource_table.scala 367:41 372:33]
  wire [30:0] _GEN_129 = rem_entry_is_last ? _GEN_95 : _res_table_wr_reg_T_24; // @[resource_table.scala 367:41 373:34]
  wire [1:0] _GEN_131 = rem_entry_is_first ? _GEN_93 : _GEN_127; // @[resource_table.scala 364:37]
  wire  _GEN_132 = rem_entry_is_first ? _GEN_94 : _GEN_128; // @[resource_table.scala 364:37]
  wire [30:0] _GEN_133 = rem_entry_is_first ? _GEN_95 : _GEN_129; // @[resource_table.scala 364:37]
  wire [30:0] _res_table_wr_reg_T_28 = {res_table_rd_reg[30:29],2'h2,rtrr_res_size,rtrr_res_strt}; // @[Cat.scala 31:58]
  wire [30:0] _res_table_wr_reg_T_32 = {2'h3,res_table_rd_reg[28:27],rtrr_res_size,rtrr_res_strt}; // @[Cat.scala 31:58]
  wire [30:0] _res_table_wr_reg_T_36 = {res_table_rd_reg[30:29],res_addr_wg_slot,rtrr_res_size,rtrr_res_strt}; // @[Cat.scala 31:58]
  wire [30:0] _GEN_135 = rem_entry_is_last ? _res_table_wr_reg_T_32 : _res_table_wr_reg_T_36; // @[resource_table.scala 385:41 389:34 393:34]
  wire [1:0] _GEN_136 = rem_entry_is_last ? _GEN_93 : res_table_wr_reg[30:29]; // @[resource_table.scala 385:41 392:34]
  wire [1:0] _GEN_137 = rem_entry_is_first ? res_addr_wg_slot : _GEN_96; // @[resource_table.scala 381:37 382:38]
  wire [30:0] _GEN_138 = rem_entry_is_first ? _res_table_wr_reg_T_28 : _GEN_135; // @[resource_table.scala 381:37 383:34]
  wire [1:0] _GEN_140 = rem_entry_is_first ? _GEN_93 : _GEN_136; // @[resource_table.scala 381:37]
  wire [1:0] _GEN_142 = 5'h10 == d_state ? _GEN_137 : _GEN_96; // @[resource_table.scala 315:20]
  wire [30:0] _GEN_143 = 5'h10 == d_state ? _GEN_138 : _GEN_95; // @[resource_table.scala 315:20]
  wire [1:0] _GEN_144 = 5'h10 == d_state ? _GEN_140 : _GEN_93; // @[resource_table.scala 315:20]
  wire [4:0] _GEN_146 = 5'h10 == d_state ? 5'h1 : d_state; // @[resource_table.scala 315:20 396:21 118:26]
  wire [4:0] _GEN_147 = 5'h8 == d_state ? 5'h10 : _GEN_146; // @[resource_table.scala 315:20]
  wire [1:0] _GEN_148 = 5'h8 == d_state ? _GEN_131 : _GEN_144; // @[resource_table.scala 315:20]
  wire  _GEN_149 = 5'h8 == d_state ? _GEN_132 : 5'h10 == d_state | _GEN_94; // @[resource_table.scala 315:20]
  wire [30:0] _GEN_150 = 5'h8 == d_state ? _GEN_133 : _GEN_143; // @[resource_table.scala 315:20]
  wire [1:0] _GEN_151 = 5'h8 == d_state ? _GEN_96 : _GEN_142; // @[resource_table.scala 315:20]
  wire  _GEN_152 = 5'h8 == d_state ? 1'h0 : 5'h10 == d_state; // @[resource_table.scala 314:18 315:20]
  wire  _GEN_153 = 5'h4 == d_state | _GEN_92; // @[resource_table.scala 315:20 355:29]
  wire [1:0] _GEN_154 = 5'h4 == d_state ? res_table_rd_reg[30:29] : _GEN_148; // @[resource_table.scala 315:20 356:30]
  wire [1:0] _GEN_158 = 5'h4 == d_state ? _GEN_96 : _GEN_151; // @[resource_table.scala 315:20]
  wire  _GEN_165 = 5'h2 == d_state ? _GEN_124 : _GEN_153; // @[resource_table.scala 315:20]
  wire [1:0] _GEN_166 = 5'h2 == d_state ? _GEN_125 : _GEN_154; // @[resource_table.scala 315:20]
  wire  _GEN_171 = 5'h1 == d_state ? _GEN_100 : _GEN_165; // @[resource_table.scala 315:20]
  wire [1:0] _GEN_172 = 5'h1 == d_state ? _GEN_101 : _GEN_166; // @[resource_table.scala 315:20]
  wire [12:0] _GEN_179 = _T_5 ? 13'h1000 : 13'h0; // @[resource_table.scala 406:36 408:69 410:40]
  wire [12:0] _GEN_180 = _T_5 ? 13'h0 : res_table_max_start; // @[resource_table.scala 138:38 408:69 411:41]
  wire  _GEN_185 = find_max_start & _T_5; // @[resource_table.scala 401:19 404:33]
  wire [12:0] _GEN_186 = find_max_start ? _GEN_180 : res_table_max_start; // @[resource_table.scala 404:33 138:38]
  wire  _T_36 = res_table_rd_reg[30:29] != 2'h3; // @[resource_table.scala 430:62]
  wire  _GEN_190 = res_table_rd_reg[30:29] != 2'h3 | _GEN_171; // @[resource_table.scala 430:88 431:37]
  wire [1:0] _GEN_191 = res_table_rd_reg[30:29] != 2'h3 ? res_table_rd_reg[30:29] : _GEN_172; // @[resource_table.scala 430:88 432:38]
  wire [3:0] _GEN_192 = res_table_rd_reg[30:29] != 2'h3 ? 4'h4 : 4'h8; // @[resource_table.scala 430:88 433:29 436:29]
  wire [12:0] _GEN_194 = res_table_rd_valid ? 13'h0 : res_table_max_start; // @[resource_table.scala 426:37 428:37 138:38]
  wire  _GEN_195 = res_table_rd_valid ? _GEN_190 : _GEN_171; // @[resource_table.scala 426:37]
  wire [1:0] _GEN_196 = res_table_rd_valid ? _GEN_191 : _GEN_172; // @[resource_table.scala 426:37]
  wire [3:0] _GEN_200 = _T_36 ? f_state : 4'h8; // @[resource_table.scala 126:26 443:88 448:29]
  wire [13:0] _GEN_292 = {{1'd0}, rtlrr_res_strt}; // @[resource_table.scala 70:89]
  wire [13:0] _T_44 = _GEN_292 + rtlrr_res_size; // @[resource_table.scala 70:89]
  wire [13:0] _GEN_293 = {{1'd0}, rtrr_res_strt}; // @[resource_table.scala 70:45]
  wire [13:0] _T_46 = _GEN_293 - _T_44; // @[resource_table.scala 70:45]
  wire [13:0] _GEN_201 = _T_46 > res_table_max_size ? _T_46 : res_table_max_size; // @[resource_table.scala 451:102 137:37 452:40]
  wire [13:0] _GEN_202 = _T_46 > res_table_max_size ? _T_44 : {{1'd0}, res_table_max_start}; // @[resource_table.scala 451:102 138:38 453:41]
  wire [3:0] _GEN_205 = res_table_rd_valid ? _GEN_200 : f_state; // @[resource_table.scala 126:26 441:37]
  wire [13:0] _GEN_206 = res_table_rd_valid ? _GEN_201 : res_table_max_size; // @[resource_table.scala 137:37 441:37]
  wire [13:0] _GEN_207 = res_table_rd_valid ? _GEN_202 : {{1'd0}, res_table_max_start}; // @[resource_table.scala 441:37 138:38]
  wire [13:0] _T_52 = _GEN_293 + rtrr_res_size; // @[resource_table.scala 73:67]
  wire [13:0] _T_54 = 14'h1000 - _T_52; // @[resource_table.scala 73:28]
  wire [13:0] _GEN_208 = _T_54 > res_table_max_size ? _T_54 : res_table_max_size; // @[resource_table.scala 459:80 460:36 137:37]
  wire [13:0] _GEN_209 = _T_54 > res_table_max_size ? _T_52 : {{1'd0}, res_table_max_start}; // @[resource_table.scala 459:80 461:37 138:38]
  wire [13:0] _GEN_210 = 4'h8 == f_state ? _GEN_208 : res_table_max_size; // @[resource_table.scala 402:20 137:37]
  wire [13:0] _GEN_211 = 4'h8 == f_state ? _GEN_209 : {{1'd0}, res_table_max_start}; // @[resource_table.scala 402:20 138:38]
  wire [3:0] _GEN_213 = 4'h8 == f_state ? 4'h1 : f_state; // @[resource_table.scala 402:20 464:21 126:26]
  wire [13:0] _GEN_218 = 4'h4 == f_state ? _GEN_207 : _GEN_211; // @[resource_table.scala 402:20]
  wire [13:0] _GEN_221 = 4'h2 == f_state ? {{1'd0}, _GEN_194} : _GEN_218; // @[resource_table.scala 402:20]
  wire [13:0] _GEN_228 = 4'h1 == f_state ? {{1'd0}, _GEN_186} : _GEN_221; // @[resource_table.scala 402:20]
  wire  _GEN_238 = ~res_addr_cu_id | cu_initialized_0; // @[resource_table.scala 151:33 476:{40,40}]
  wire  _GEN_239 = res_addr_cu_id | cu_initialized_1; // @[resource_table.scala 151:33 476:{40,40}]
  wire [3:0] _res_table_rd_reg_T = 3'h4 * res_addr_cu_id; // @[resource_table.scala 50:34]
  wire [3:0] _GEN_301 = {{2'd0}, res_addr_wg_slot}; // @[resource_table.scala 50:42]
  wire [3:0] _res_table_rd_reg_T_2 = _res_table_rd_reg_T + _GEN_301; // @[resource_table.scala 50:42]
  wire [30:0] _GEN_251 = 4'h1 == _res_table_rd_reg_T_2 ? resource_table_ram_1 : resource_table_ram_0; // @[resource_table.scala 480:{26,26}]
  wire [30:0] _GEN_252 = 4'h2 == _res_table_rd_reg_T_2 ? resource_table_ram_2 : _GEN_251; // @[resource_table.scala 480:{26,26}]
  wire [30:0] _GEN_253 = 4'h3 == _res_table_rd_reg_T_2 ? resource_table_ram_3 : _GEN_252; // @[resource_table.scala 480:{26,26}]
  wire [30:0] _GEN_254 = 4'h4 == _res_table_rd_reg_T_2 ? resource_table_ram_4 : _GEN_253; // @[resource_table.scala 480:{26,26}]
  wire [30:0] _GEN_255 = 4'h5 == _res_table_rd_reg_T_2 ? resource_table_ram_5 : _GEN_254; // @[resource_table.scala 480:{26,26}]
  wire [30:0] _GEN_256 = 4'h6 == _res_table_rd_reg_T_2 ? resource_table_ram_6 : _GEN_255; // @[resource_table.scala 480:{26,26}]
  wire [30:0] _GEN_257 = 4'h7 == _res_table_rd_reg_T_2 ? resource_table_ram_7 : _GEN_256; // @[resource_table.scala 480:{26,26}]
  wire [13:0] _GEN_303 = reset ? 14'h0 : _GEN_228; // @[resource_table.scala 138:{38,38}]
  assign io_res_table_done_o = res_table_done; // @[resource_table.scala 25:25]
  assign io_cam_biggest_space_size = res_table_max_size; // @[resource_table.scala 486:31]
  assign io_cam_biggest_space_addr = res_table_max_start; // @[resource_table.scala 487:31]
  always @(posedge clock) begin
    if (reset) begin // @[resource_table.scala 24:33]
      res_table_done <= 1'h0; // @[resource_table.scala 24:33]
    end else if (4'h1 == m_state) begin // @[resource_table.scala 190:20]
      res_table_done <= 1'h0; // @[resource_table.scala 189:20]
    end else if (4'h2 == m_state) begin // @[resource_table.scala 190:20]
      res_table_done <= 1'h0; // @[resource_table.scala 189:20]
    end else if (4'h4 == m_state) begin // @[resource_table.scala 190:20]
      res_table_done <= 1'h0; // @[resource_table.scala 189:20]
    end else begin
      res_table_done <= 4'h8 == m_state & find_max_done;
    end
    if (reset) begin // @[resource_table.scala 39:33]
      alloc_res_en_i <= 1'h0; // @[resource_table.scala 39:33]
    end else begin
      alloc_res_en_i <= io_alloc_res_en; // @[resource_table.scala 169:20]
    end
    if (reset) begin // @[resource_table.scala 40:35]
      dealloc_res_en_i <= 1'h0; // @[resource_table.scala 40:35]
    end else begin
      dealloc_res_en_i <= io_dealloc_res_en; // @[resource_table.scala 178:22]
    end
    if (reset) begin // @[resource_table.scala 43:37]
      alloc_wg_slot_id_i <= 2'h0; // @[resource_table.scala 43:37]
    end else if (io_alloc_res_en) begin // @[resource_table.scala 170:26]
      alloc_wg_slot_id_i <= io_alloc_wg_slot_id; // @[resource_table.scala 172:28]
    end
    if (reset) begin // @[resource_table.scala 44:39]
      dealloc_wg_slot_id_i <= 2'h0; // @[resource_table.scala 44:39]
    end else if (io_dealloc_res_en) begin // @[resource_table.scala 179:28]
      dealloc_wg_slot_id_i <= io_dealloc_wg_slot_id; // @[resource_table.scala 181:30]
    end
    if (reset) begin // @[resource_table.scala 46:35]
      alloc_res_size_i <= 14'h0; // @[resource_table.scala 46:35]
    end else if (io_alloc_res_en) begin // @[resource_table.scala 170:26]
      alloc_res_size_i <= io_alloc_res_size; // @[resource_table.scala 173:26]
    end
    if (reset) begin // @[resource_table.scala 47:36]
      alloc_res_start_i <= 13'h0; // @[resource_table.scala 47:36]
    end else if (io_alloc_res_en) begin // @[resource_table.scala 170:26]
      alloc_res_start_i <= io_alloc_res_start; // @[resource_table.scala 174:27]
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_0 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h0 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_0 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_1 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h1 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_1 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_2 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h2 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_2 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_3 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h3 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_3 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_4 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h4 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_4 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_5 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h5 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_5 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_6 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h6 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_6 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_7 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h7 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_7 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_8 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h8 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_8 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 80:37]
      resource_table_ram_9 <= 31'h0; // @[resource_table.scala 80:37]
    end else if (!(res_table_rd_en)) begin // @[resource_table.scala 479:26]
      if (res_table_wr_en) begin // @[resource_table.scala 483:31]
        if (4'h9 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 484:79]
          resource_table_ram_9 <= res_table_wr_reg; // @[resource_table.scala 484:79]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 81:37]
      table_head_pointer_0 <= 2'h0; // @[resource_table.scala 81:37]
    end else if (!(alloc_res_en_i | dealloc_res_en_i)) begin // @[resource_table.scala 468:45]
      if (alloc_done | dealloc_done) begin // @[resource_table.scala 473:42]
        if (~res_addr_cu_id) begin // @[resource_table.scala 475:44]
          table_head_pointer_0 <= table_head_pointer_i; // @[resource_table.scala 475:44]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 81:37]
      table_head_pointer_1 <= 2'h0; // @[resource_table.scala 81:37]
    end else if (!(alloc_res_en_i | dealloc_res_en_i)) begin // @[resource_table.scala 468:45]
      if (alloc_done | dealloc_done) begin // @[resource_table.scala 473:42]
        if (res_addr_cu_id) begin // @[resource_table.scala 475:44]
          table_head_pointer_1 <= table_head_pointer_i; // @[resource_table.scala 475:44]
        end
      end
    end
    if (reset) begin // @[resource_table.scala 82:39]
      table_head_pointer_i <= 2'h0; // @[resource_table.scala 82:39]
    end else if (alloc_res_en_i | dealloc_res_en_i) begin // @[resource_table.scala 468:45]
      if (res_addr_cu_id) begin // @[resource_table.scala 471:30]
        table_head_pointer_i <= table_head_pointer_1; // @[resource_table.scala 471:30]
      end else begin
        table_head_pointer_i <= table_head_pointer_0;
      end
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      if (!(4'h1 == a_state)) begin // @[resource_table.scala 228:20]
        table_head_pointer_i <= _GEN_87;
      end
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      table_head_pointer_i <= _GEN_119;
    end else begin
      table_head_pointer_i <= _GEN_158;
    end
    if (reset) begin // @[resource_table.scala 103:26]
      m_state <= 4'h1; // @[resource_table.scala 103:26]
    end else if (4'h1 == m_state) begin // @[resource_table.scala 190:20]
      if (alloc_res_en_i) begin // @[resource_table.scala 192:33]
        m_state <= 4'h2; // @[resource_table.scala 194:25]
      end else if (dealloc_res_en_i) begin // @[resource_table.scala 196:40]
        m_state <= 4'h4; // @[resource_table.scala 198:25]
      end
    end else if (4'h2 == m_state) begin // @[resource_table.scala 190:20]
      if (alloc_done) begin // @[resource_table.scala 202:29]
        m_state <= 4'h8; // @[resource_table.scala 204:25]
      end
    end else if (4'h4 == m_state) begin // @[resource_table.scala 190:20]
      m_state <= _GEN_16;
    end else begin
      m_state <= _GEN_20;
    end
    if (reset) begin // @[resource_table.scala 110:26]
      a_state <= 4'h1; // @[resource_table.scala 110:26]
    end else if (4'h1 == a_state) begin // @[resource_table.scala 228:20]
      if (alloc_start) begin // @[resource_table.scala 230:30]
        if (table_head_pointer_i == 2'h3 | ~cu_initialized_i) begin // @[resource_table.scala 235:90]
          a_state <= 4'h8; // @[resource_table.scala 238:29]
        end else begin
          a_state <= 4'h2; // @[resource_table.scala 245:29]
        end
      end
    end else if (4'h2 == a_state) begin // @[resource_table.scala 228:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 251:37]
        a_state <= _GEN_54;
      end
    end else if (4'h4 == a_state) begin // @[resource_table.scala 228:20]
      a_state <= 4'h8; // @[resource_table.scala 286:21]
    end else begin
      a_state <= _GEN_73;
    end
    if (reset) begin // @[resource_table.scala 118:26]
      d_state <= 5'h1; // @[resource_table.scala 118:26]
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      if (dealloc_start) begin // @[resource_table.scala 317:32]
        d_state <= 5'h2; // @[resource_table.scala 322:25]
      end
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 327:37]
        d_state <= {{1'd0}, _GEN_114};
      end
    end else if (5'h4 == d_state) begin // @[resource_table.scala 315:20]
      d_state <= 5'h8; // @[resource_table.scala 357:21]
    end else begin
      d_state <= _GEN_147;
    end
    if (reset) begin // @[resource_table.scala 126:26]
      f_state <= 4'h1; // @[resource_table.scala 126:26]
    end else if (4'h1 == f_state) begin // @[resource_table.scala 402:20]
      if (find_max_start) begin // @[resource_table.scala 404:33]
        if (!(_T_5)) begin // @[resource_table.scala 408:69]
          f_state <= 4'h2; // @[resource_table.scala 417:29]
        end
      end
    end else if (4'h2 == f_state) begin // @[resource_table.scala 402:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 426:37]
        f_state <= _GEN_192;
      end
    end else if (4'h4 == f_state) begin // @[resource_table.scala 402:20]
      f_state <= _GEN_205;
    end else begin
      f_state <= _GEN_213;
    end
    if (reset) begin // @[resource_table.scala 129:35]
      res_table_wr_reg <= 31'h0; // @[resource_table.scala 129:35]
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      res_table_wr_reg <= _GEN_95;
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      res_table_wr_reg <= _GEN_95;
    end else if (5'h4 == d_state) begin // @[resource_table.scala 315:20]
      res_table_wr_reg <= _GEN_95;
    end else begin
      res_table_wr_reg <= _GEN_150;
    end
    if (reset) begin // @[resource_table.scala 130:35]
      res_table_rd_reg <= 31'h0; // @[resource_table.scala 130:35]
    end else if (res_table_rd_en) begin // @[resource_table.scala 479:26]
      if (4'h9 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 480:26]
        res_table_rd_reg <= resource_table_ram_9; // @[resource_table.scala 480:26]
      end else if (4'h8 == _res_table_rd_reg_T_2) begin // @[resource_table.scala 480:26]
        res_table_rd_reg <= resource_table_ram_8; // @[resource_table.scala 480:26]
      end else begin
        res_table_rd_reg <= _GEN_257;
      end
    end
    if (reset) begin // @[resource_table.scala 131:40]
      res_table_last_rd_reg <= 31'h0; // @[resource_table.scala 131:40]
    end else if (res_table_rd_en) begin // @[resource_table.scala 479:26]
      res_table_last_rd_reg <= res_table_rd_reg; // @[resource_table.scala 481:31]
    end
    if (reset) begin // @[resource_table.scala 132:33]
      res_addr_cu_id <= 1'h0; // @[resource_table.scala 132:33]
    end else if (io_dealloc_res_en) begin // @[resource_table.scala 179:28]
      res_addr_cu_id <= io_dealloc_cu_id; // @[resource_table.scala 182:24]
    end else if (io_alloc_res_en) begin // @[resource_table.scala 170:26]
      res_addr_cu_id <= io_alloc_cu_id; // @[resource_table.scala 175:24]
    end
    if (reset) begin // @[resource_table.scala 133:35]
      res_addr_wg_slot <= 2'h0; // @[resource_table.scala 133:35]
    end else if (4'h1 == f_state) begin // @[resource_table.scala 402:20]
      if (find_max_start) begin // @[resource_table.scala 404:33]
        if (_T_5) begin // @[resource_table.scala 408:69]
          res_addr_wg_slot <= _GEN_172;
        end else begin
          res_addr_wg_slot <= table_head_pointer_i; // @[resource_table.scala 416:38]
        end
      end else begin
        res_addr_wg_slot <= _GEN_172;
      end
    end else if (4'h2 == f_state) begin // @[resource_table.scala 402:20]
      res_addr_wg_slot <= _GEN_196;
    end else if (4'h4 == f_state) begin // @[resource_table.scala 402:20]
      res_addr_wg_slot <= _GEN_196;
    end else begin
      res_addr_wg_slot <= _GEN_172;
    end
    if (reset) begin // @[resource_table.scala 134:34]
      res_table_rd_en <= 1'h0; // @[resource_table.scala 134:34]
    end else if (4'h1 == f_state) begin // @[resource_table.scala 402:20]
      if (find_max_start) begin // @[resource_table.scala 404:33]
        if (_T_5) begin // @[resource_table.scala 408:69]
          res_table_rd_en <= _GEN_171;
        end else begin
          res_table_rd_en <= 1'h1; // @[resource_table.scala 415:37]
        end
      end else begin
        res_table_rd_en <= _GEN_171;
      end
    end else if (4'h2 == f_state) begin // @[resource_table.scala 402:20]
      res_table_rd_en <= _GEN_195;
    end else if (4'h4 == f_state) begin // @[resource_table.scala 402:20]
      res_table_rd_en <= _GEN_195;
    end else begin
      res_table_rd_en <= _GEN_171;
    end
    if (reset) begin // @[resource_table.scala 135:34]
      res_table_wr_en <= 1'h0; // @[resource_table.scala 135:34]
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      res_table_wr_en <= _GEN_94;
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      res_table_wr_en <= _GEN_94;
    end else if (5'h4 == d_state) begin // @[resource_table.scala 315:20]
      res_table_wr_en <= _GEN_94;
    end else begin
      res_table_wr_en <= _GEN_149;
    end
    if (reset) begin // @[resource_table.scala 136:37]
      res_table_rd_valid <= 1'h0; // @[resource_table.scala 136:37]
    end else begin
      res_table_rd_valid <= res_table_rd_en; // @[resource_table.scala 478:24]
    end
    if (reset) begin // @[resource_table.scala 137:37]
      res_table_max_size <= 14'h0; // @[resource_table.scala 137:37]
    end else if (4'h1 == f_state) begin // @[resource_table.scala 402:20]
      if (find_max_start) begin // @[resource_table.scala 404:33]
        res_table_max_size <= {{1'd0}, _GEN_179};
      end
    end else if (4'h2 == f_state) begin // @[resource_table.scala 402:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 426:37]
        res_table_max_size <= {{1'd0}, rtrr_res_strt}; // @[resource_table.scala 427:36]
      end
    end else if (4'h4 == f_state) begin // @[resource_table.scala 402:20]
      res_table_max_size <= _GEN_206;
    end else begin
      res_table_max_size <= _GEN_210;
    end
    res_table_max_start <= _GEN_303[12:0]; // @[resource_table.scala 138:{38,38}]
    if (reset) begin // @[resource_table.scala 141:30]
      alloc_start <= 1'h0; // @[resource_table.scala 141:30]
    end else begin
      alloc_start <= _GEN_27;
    end
    if (reset) begin // @[resource_table.scala 142:32]
      dealloc_start <= 1'h0; // @[resource_table.scala 142:32]
    end else begin
      dealloc_start <= _GEN_29;
    end
    if (reset) begin // @[resource_table.scala 143:33]
      find_max_start <= 1'h0; // @[resource_table.scala 143:33]
    end else if (4'h1 == m_state) begin // @[resource_table.scala 190:20]
      find_max_start <= 1'h0; // @[resource_table.scala 188:20]
    end else if (4'h2 == m_state) begin // @[resource_table.scala 190:20]
      find_max_start <= alloc_done;
    end else begin
      find_max_start <= _GEN_21;
    end
    if (reset) begin // @[resource_table.scala 144:29]
      alloc_done <= 1'h0; // @[resource_table.scala 144:29]
    end else if (4'h1 == a_state) begin // @[resource_table.scala 228:20]
      alloc_done <= 1'h0; // @[resource_table.scala 226:16]
    end else if (4'h2 == a_state) begin // @[resource_table.scala 228:20]
      alloc_done <= 1'h0; // @[resource_table.scala 226:16]
    end else if (4'h4 == a_state) begin // @[resource_table.scala 228:20]
      alloc_done <= 1'h0; // @[resource_table.scala 226:16]
    end else begin
      alloc_done <= 4'h8 == a_state;
    end
    if (reset) begin // @[resource_table.scala 145:31]
      dealloc_done <= 1'h0; // @[resource_table.scala 145:31]
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      dealloc_done <= 1'h0; // @[resource_table.scala 314:18]
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      dealloc_done <= _GEN_120;
    end else if (5'h4 == d_state) begin // @[resource_table.scala 315:20]
      dealloc_done <= 1'h0; // @[resource_table.scala 314:18]
    end else begin
      dealloc_done <= _GEN_152;
    end
    if (reset) begin // @[resource_table.scala 146:32]
      find_max_done <= 1'h0; // @[resource_table.scala 146:32]
    end else if (4'h1 == f_state) begin // @[resource_table.scala 402:20]
      find_max_done <= _GEN_185;
    end else if (4'h2 == f_state) begin // @[resource_table.scala 402:20]
      find_max_done <= 1'h0; // @[resource_table.scala 401:19]
    end else if (4'h4 == f_state) begin // @[resource_table.scala 402:20]
      find_max_done <= 1'h0; // @[resource_table.scala 401:19]
    end else begin
      find_max_done <= 4'h8 == f_state;
    end
    if (reset) begin // @[resource_table.scala 147:36]
      new_entry_is_last <= 1'h0; // @[resource_table.scala 147:36]
    end else if (4'h1 == a_state) begin // @[resource_table.scala 228:20]
      if (alloc_start) begin // @[resource_table.scala 230:30]
        new_entry_is_last <= _T_7;
      end
    end else if (4'h2 == a_state) begin // @[resource_table.scala 228:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 251:37]
        new_entry_is_last <= _GEN_55;
      end
    end
    if (reset) begin // @[resource_table.scala 148:37]
      new_entry_is_first <= 1'h0; // @[resource_table.scala 148:37]
    end else if (4'h1 == a_state) begin // @[resource_table.scala 228:20]
      if (alloc_start) begin // @[resource_table.scala 230:30]
        new_entry_is_first <= _T_7;
      end
    end else if (4'h2 == a_state) begin // @[resource_table.scala 228:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 251:37]
        new_entry_is_first <= _GEN_51;
      end
    end
    if (reset) begin // @[resource_table.scala 149:36]
      rem_entry_is_last <= 1'h0; // @[resource_table.scala 149:36]
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      if (dealloc_start) begin // @[resource_table.scala 317:32]
        rem_entry_is_last <= 1'h0; // @[resource_table.scala 319:35]
      end
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 327:37]
        rem_entry_is_last <= _GEN_116;
      end
    end
    if (reset) begin // @[resource_table.scala 150:37]
      rem_entry_is_first <= 1'h0; // @[resource_table.scala 150:37]
    end else if (5'h1 == d_state) begin // @[resource_table.scala 315:20]
      if (dealloc_start) begin // @[resource_table.scala 317:32]
        rem_entry_is_first <= 1'h0; // @[resource_table.scala 318:36]
      end
    end else if (5'h2 == d_state) begin // @[resource_table.scala 315:20]
      if (res_table_rd_valid) begin // @[resource_table.scala 327:37]
        rem_entry_is_first <= _GEN_115;
      end
    end
    if (reset) begin // @[resource_table.scala 151:33]
      cu_initialized_0 <= 1'h0; // @[resource_table.scala 151:33]
    end else if (!(alloc_res_en_i | dealloc_res_en_i)) begin // @[resource_table.scala 468:45]
      if (alloc_done | dealloc_done) begin // @[resource_table.scala 473:42]
        cu_initialized_0 <= _GEN_238;
      end
    end
    if (reset) begin // @[resource_table.scala 151:33]
      cu_initialized_1 <= 1'h0; // @[resource_table.scala 151:33]
    end else if (!(alloc_res_en_i | dealloc_res_en_i)) begin // @[resource_table.scala 468:45]
      if (alloc_done | dealloc_done) begin // @[resource_table.scala 473:42]
        cu_initialized_1 <= _GEN_239;
      end
    end
    if (reset) begin // @[resource_table.scala 152:35]
      cu_initialized_i <= 1'h0; // @[resource_table.scala 152:35]
    end else if (alloc_res_en_i | dealloc_res_en_i) begin // @[resource_table.scala 468:45]
      if (res_addr_cu_id) begin // @[resource_table.scala 470:26]
        cu_initialized_i <= cu_initialized_1; // @[resource_table.scala 470:26]
      end else begin
        cu_initialized_i <= cu_initialized_0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  res_table_done = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  alloc_res_en_i = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  dealloc_res_en_i = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alloc_wg_slot_id_i = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  dealloc_wg_slot_id_i = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  alloc_res_size_i = _RAND_5[13:0];
  _RAND_6 = {1{`RANDOM}};
  alloc_res_start_i = _RAND_6[12:0];
  _RAND_7 = {1{`RANDOM}};
  resource_table_ram_0 = _RAND_7[30:0];
  _RAND_8 = {1{`RANDOM}};
  resource_table_ram_1 = _RAND_8[30:0];
  _RAND_9 = {1{`RANDOM}};
  resource_table_ram_2 = _RAND_9[30:0];
  _RAND_10 = {1{`RANDOM}};
  resource_table_ram_3 = _RAND_10[30:0];
  _RAND_11 = {1{`RANDOM}};
  resource_table_ram_4 = _RAND_11[30:0];
  _RAND_12 = {1{`RANDOM}};
  resource_table_ram_5 = _RAND_12[30:0];
  _RAND_13 = {1{`RANDOM}};
  resource_table_ram_6 = _RAND_13[30:0];
  _RAND_14 = {1{`RANDOM}};
  resource_table_ram_7 = _RAND_14[30:0];
  _RAND_15 = {1{`RANDOM}};
  resource_table_ram_8 = _RAND_15[30:0];
  _RAND_16 = {1{`RANDOM}};
  resource_table_ram_9 = _RAND_16[30:0];
  _RAND_17 = {1{`RANDOM}};
  table_head_pointer_0 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  table_head_pointer_1 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  table_head_pointer_i = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  m_state = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  a_state = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  d_state = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  f_state = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  res_table_wr_reg = _RAND_24[30:0];
  _RAND_25 = {1{`RANDOM}};
  res_table_rd_reg = _RAND_25[30:0];
  _RAND_26 = {1{`RANDOM}};
  res_table_last_rd_reg = _RAND_26[30:0];
  _RAND_27 = {1{`RANDOM}};
  res_addr_cu_id = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  res_addr_wg_slot = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  res_table_rd_en = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  res_table_wr_en = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  res_table_rd_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  res_table_max_size = _RAND_32[13:0];
  _RAND_33 = {1{`RANDOM}};
  res_table_max_start = _RAND_33[12:0];
  _RAND_34 = {1{`RANDOM}};
  alloc_start = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dealloc_start = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  find_max_start = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  alloc_done = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dealloc_done = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  find_max_done = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  new_entry_is_last = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  new_entry_is_first = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  rem_entry_is_last = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  rem_entry_is_first = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  cu_initialized_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  cu_initialized_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  cu_initialized_i = _RAND_46[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module wg_resource_table_neo(
  input        clock,
  input        reset,
  output [2:0] io_wf_count_out,
  input        io_cu_id,
  input        io_alloc_en,
  input        io_dealloc_en,
  input  [2:0] io_wf_count_in,
  input  [1:0] io_alloc_wg_slot_id,
  input  [1:0] io_dealloc_wg_slot_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] wf_count_out_i_0; // @[wg_resource_table_neo.scala 15:33]
  reg [2:0] wf_count_out_i_1; // @[wg_resource_table_neo.scala 15:33]
  reg [2:0] wf_count_per_wg_slot_0_0; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_0_1; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_0_2; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_0_3; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_1_0; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_1_1; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_1_2; // @[wg_resource_table_neo.scala 16:39]
  reg [2:0] wf_count_per_wg_slot_1_3; // @[wg_resource_table_neo.scala 16:39]
  wire [2:0] _GEN_1 = io_cu_id ? wf_count_out_i_1 : wf_count_out_i_0; // @[wg_resource_table_neo.scala 26:{62,62}]
  wire [2:0] _wf_count_out_i_T_1 = _GEN_1 - io_wf_count_in; // @[wg_resource_table_neo.scala 26:62]
  wire  _GEN_36 = ~io_cu_id; // @[wg_resource_table_neo.scala 16:39 27:{61,61}]
  wire [2:0] _GEN_13 = _GEN_36 & 2'h1 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_0_1 : wf_count_per_wg_slot_0_0; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _GEN_14 = _GEN_36 & 2'h2 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_0_2 : _GEN_13; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _GEN_15 = _GEN_36 & 2'h3 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_0_3 : _GEN_14; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _GEN_16 = io_cu_id & 2'h0 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_1_0 : _GEN_15; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _GEN_17 = io_cu_id & 2'h1 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_1_1 : _GEN_16; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _GEN_18 = io_cu_id & 2'h2 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_1_2 : _GEN_17; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _GEN_19 = io_cu_id & 2'h3 == io_dealloc_wg_slot_id ? wf_count_per_wg_slot_1_3 : _GEN_18; // @[wg_resource_table_neo.scala 31:{62,62}]
  wire [2:0] _wf_count_out_i_T_3 = _GEN_1 + _GEN_19; // @[wg_resource_table_neo.scala 31:62]
  reg  cu_id_delay; // @[wg_resource_table_neo.scala 34:30]
  assign io_wf_count_out = cu_id_delay ? wf_count_out_i_1 : wf_count_out_i_0; // @[wg_resource_table_neo.scala 36:{21,21}]
  always @(posedge clock) begin
    if (reset) begin // @[wg_resource_table_neo.scala 15:33]
      wf_count_out_i_0 <= 3'h4; // @[wg_resource_table_neo.scala 15:33]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (~io_cu_id) begin // @[wg_resource_table_neo.scala 26:34]
        wf_count_out_i_0 <= _wf_count_out_i_T_1; // @[wg_resource_table_neo.scala 26:34]
      end
    end else if (io_dealloc_en) begin // @[wg_resource_table_neo.scala 30:29]
      if (~io_cu_id) begin // @[wg_resource_table_neo.scala 31:34]
        wf_count_out_i_0 <= _wf_count_out_i_T_3; // @[wg_resource_table_neo.scala 31:34]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 15:33]
      wf_count_out_i_1 <= 3'h4; // @[wg_resource_table_neo.scala 15:33]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (io_cu_id) begin // @[wg_resource_table_neo.scala 26:34]
        wf_count_out_i_1 <= _wf_count_out_i_T_1; // @[wg_resource_table_neo.scala 26:34]
      end
    end else if (io_dealloc_en) begin // @[wg_resource_table_neo.scala 30:29]
      if (io_cu_id) begin // @[wg_resource_table_neo.scala 31:34]
        wf_count_out_i_1 <= _wf_count_out_i_T_3; // @[wg_resource_table_neo.scala 31:34]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_0_0 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (~io_cu_id & 2'h0 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_0_0 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_0_1 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (~io_cu_id & 2'h1 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_0_1 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_0_2 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (~io_cu_id & 2'h2 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_0_2 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_0_3 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (~io_cu_id & 2'h3 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_0_3 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_1_0 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (io_cu_id & 2'h0 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_1_0 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_1_1 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (io_cu_id & 2'h1 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_1_1 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_1_2 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (io_cu_id & 2'h2 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_1_2 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 16:39]
      wf_count_per_wg_slot_1_3 <= 3'h0; // @[wg_resource_table_neo.scala 16:39]
    end else if (io_alloc_en) begin // @[wg_resource_table_neo.scala 25:22]
      if (io_cu_id & 2'h3 == io_alloc_wg_slot_id) begin // @[wg_resource_table_neo.scala 27:61]
        wf_count_per_wg_slot_1_3 <= io_wf_count_in; // @[wg_resource_table_neo.scala 27:61]
      end
    end
    if (reset) begin // @[wg_resource_table_neo.scala 34:30]
      cu_id_delay <= 1'h0; // @[wg_resource_table_neo.scala 34:30]
    end else begin
      cu_id_delay <= io_cu_id; // @[wg_resource_table_neo.scala 35:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wf_count_out_i_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  wf_count_out_i_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  wf_count_per_wg_slot_0_0 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  wf_count_per_wg_slot_0_1 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  wf_count_per_wg_slot_0_2 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  wf_count_per_wg_slot_0_3 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  wf_count_per_wg_slot_1_0 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  wf_count_per_wg_slot_1_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  wf_count_per_wg_slot_1_2 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  wf_count_per_wg_slot_1_3 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  cu_id_delay = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module wg_slot_id_convert_opt(
  input        clock,
  input        reset,
  input  [4:0] io_wg_id,
  input        io_cu_id,
  output [1:0] io_wg_slot_id_gen,
  output [1:0] io_wg_slot_id_find,
  input        io_find_and_cancel,
  input        io_generate
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] wg_slot_id_find_i; // @[wg_slot_id_convert_opt.scala 15:36]
  reg [1:0] wg_slot_id_gen_i; // @[wg_slot_id_convert_opt.scala 18:35]
  reg  wg_slot_id_bitmap_0_0; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_0_1; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_0_2; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_0_3; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_1_0; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_1_1; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_1_2; // @[wg_slot_id_convert_opt.scala 20:36]
  reg  wg_slot_id_bitmap_1_3; // @[wg_slot_id_convert_opt.scala 20:36]
  wire  _GEN_1 = io_cu_id ? wg_slot_id_bitmap_1_3 : wg_slot_id_bitmap_0_3; // @[wg_slot_id_convert_opt.scala 34:{14,14}]
  wire [1:0] _GEN_2 = ~_GEN_1 ? 2'h3 : 2'h0; // @[wg_slot_id_convert_opt.scala 32:19 34:46 35:27]
  wire  _GEN_5 = io_cu_id ? wg_slot_id_bitmap_1_2 : wg_slot_id_bitmap_0_2; // @[wg_slot_id_convert_opt.scala 34:{14,14}]
  wire [1:0] _GEN_6 = ~_GEN_5 ? 2'h2 : _GEN_2; // @[wg_slot_id_convert_opt.scala 34:46 35:27]
  wire  _GEN_9 = io_cu_id ? wg_slot_id_bitmap_1_1 : wg_slot_id_bitmap_0_1; // @[wg_slot_id_convert_opt.scala 34:{14,14}]
  wire [1:0] _GEN_10 = ~_GEN_9 ? 2'h1 : _GEN_6; // @[wg_slot_id_convert_opt.scala 34:46 35:27]
  wire  _GEN_13 = io_cu_id ? wg_slot_id_bitmap_1_0 : wg_slot_id_bitmap_0_0; // @[wg_slot_id_convert_opt.scala 34:{14,14}]
  wire [1:0] first_slot_id = ~_GEN_13 ? 2'h0 : _GEN_10; // @[wg_slot_id_convert_opt.scala 34:46 35:27]
  wire  first_slot_id_valid = ~_GEN_13 | (~_GEN_9 | (~_GEN_5 | ~_GEN_1)); // @[wg_slot_id_convert_opt.scala 34:46 36:33]
  wire  _T_4 = io_generate & first_slot_id_valid; // @[wg_slot_id_convert_opt.scala 40:22]
  wire  _GEN_72 = ~io_cu_id; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_73 = 2'h0 == first_slot_id; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_16 = ~io_cu_id & 2'h0 == first_slot_id | wg_slot_id_bitmap_0_0; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_76 = 2'h1 == first_slot_id; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_17 = ~io_cu_id & 2'h1 == first_slot_id | wg_slot_id_bitmap_0_1; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_79 = 2'h2 == first_slot_id; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_18 = ~io_cu_id & 2'h2 == first_slot_id | wg_slot_id_bitmap_0_2; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_82 = 2'h3 == first_slot_id; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_19 = ~io_cu_id & 2'h3 == first_slot_id | wg_slot_id_bitmap_0_3; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_20 = io_cu_id & 2'h0 == first_slot_id | wg_slot_id_bitmap_1_0; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_21 = io_cu_id & 2'h1 == first_slot_id | wg_slot_id_bitmap_1_1; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_22 = io_cu_id & 2'h2 == first_slot_id | wg_slot_id_bitmap_1_2; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_23 = io_cu_id & 2'h3 == first_slot_id | wg_slot_id_bitmap_1_3; // @[wg_slot_id_convert_opt.scala 20:36 41:{52,52}]
  wire  _GEN_24 = io_generate & first_slot_id_valid ? _GEN_16 : wg_slot_id_bitmap_0_0; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_25 = io_generate & first_slot_id_valid ? _GEN_17 : wg_slot_id_bitmap_0_1; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_26 = io_generate & first_slot_id_valid ? _GEN_18 : wg_slot_id_bitmap_0_2; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_27 = io_generate & first_slot_id_valid ? _GEN_19 : wg_slot_id_bitmap_0_3; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_28 = io_generate & first_slot_id_valid ? _GEN_20 : wg_slot_id_bitmap_1_0; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_29 = io_generate & first_slot_id_valid ? _GEN_21 : wg_slot_id_bitmap_1_1; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_30 = io_generate & first_slot_id_valid ? _GEN_22 : wg_slot_id_bitmap_1_2; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  wire  _GEN_31 = io_generate & first_slot_id_valid ? _GEN_23 : wg_slot_id_bitmap_1_3; // @[wg_slot_id_convert_opt.scala 20:36 40:45]
  reg [4:0] wg_slot_id_find_ram_cam_0_1; // @[wg_slot_id_convert_opt.scala 52:42]
  reg [4:0] wg_slot_id_find_ram_cam_0_2; // @[wg_slot_id_convert_opt.scala 52:42]
  reg [4:0] wg_slot_id_find_ram_cam_0_3; // @[wg_slot_id_convert_opt.scala 52:42]
  reg [4:0] wg_slot_id_find_ram_cam_1_0; // @[wg_slot_id_convert_opt.scala 52:42]
  reg [4:0] wg_slot_id_find_ram_cam_1_1; // @[wg_slot_id_convert_opt.scala 52:42]
  reg [4:0] wg_slot_id_find_ram_cam_1_2; // @[wg_slot_id_convert_opt.scala 52:42]
  reg [4:0] wg_slot_id_find_ram_cam_1_3; // @[wg_slot_id_convert_opt.scala 52:42]
  wire  _T_8 = wg_slot_id_find_ram_cam_0_1 == io_wg_id & wg_slot_id_bitmap_0_1; // @[wg_slot_id_convert_opt.scala 64:61]
  wire [1:0] _GEN_34 = wg_slot_id_find_ram_cam_0_2 == io_wg_id & wg_slot_id_bitmap_0_2 ? 2'h2 : {{1'd0}, _T_8}; // @[wg_slot_id_convert_opt.scala 64:88 65:29]
  wire [1:0] _GEN_35 = wg_slot_id_find_ram_cam_0_3 == io_wg_id & wg_slot_id_bitmap_0_3 ? 2'h3 : _GEN_34; // @[wg_slot_id_convert_opt.scala 64:88 65:29]
  wire [1:0] _GEN_36 = wg_slot_id_find_ram_cam_1_0 == io_wg_id & wg_slot_id_bitmap_1_0 ? 2'h0 : _GEN_35; // @[wg_slot_id_convert_opt.scala 64:88 65:29]
  wire [1:0] _GEN_37 = wg_slot_id_find_ram_cam_1_1 == io_wg_id & wg_slot_id_bitmap_1_1 ? 2'h1 : _GEN_36; // @[wg_slot_id_convert_opt.scala 64:88 65:29]
  wire [1:0] _GEN_38 = wg_slot_id_find_ram_cam_1_2 == io_wg_id & wg_slot_id_bitmap_1_2 ? 2'h2 : _GEN_37; // @[wg_slot_id_convert_opt.scala 64:88 65:29]
  wire [1:0] _GEN_39 = wg_slot_id_find_ram_cam_1_3 == io_wg_id & wg_slot_id_bitmap_1_3 ? 2'h3 : _GEN_38; // @[wg_slot_id_convert_opt.scala 64:88 65:29]
  reg  cu_id_cancel; // @[wg_slot_id_convert_opt.scala 75:31]
  reg  cancel_valid; // @[wg_slot_id_convert_opt.scala 76:31]
  wire [4:0] found_wg_id = {{3'd0}, _GEN_39}; // @[wg_slot_id_convert_opt.scala 14:27]
  wire [4:0] _GEN_116 = reset ? 5'h0 : found_wg_id; // @[wg_slot_id_convert_opt.scala 15:{36,36} 69:23]
  assign io_wg_slot_id_gen = wg_slot_id_gen_i; // @[wg_slot_id_convert_opt.scala 19:23]
  assign io_wg_slot_id_find = wg_slot_id_find_i; // @[wg_slot_id_convert_opt.scala 16:24]
  always @(posedge clock) begin
    wg_slot_id_find_i <= _GEN_116[1:0]; // @[wg_slot_id_convert_opt.scala 15:{36,36} 69:23]
    if (reset) begin // @[wg_slot_id_convert_opt.scala 18:35]
      wg_slot_id_gen_i <= 2'h0; // @[wg_slot_id_convert_opt.scala 18:35]
    end else if (~_GEN_13) begin // @[wg_slot_id_convert_opt.scala 34:46]
      wg_slot_id_gen_i <= 2'h0; // @[wg_slot_id_convert_opt.scala 35:27]
    end else if (~_GEN_9) begin // @[wg_slot_id_convert_opt.scala 34:46]
      wg_slot_id_gen_i <= 2'h1; // @[wg_slot_id_convert_opt.scala 35:27]
    end else if (~_GEN_5) begin // @[wg_slot_id_convert_opt.scala 34:46]
      wg_slot_id_gen_i <= 2'h2; // @[wg_slot_id_convert_opt.scala 35:27]
    end else begin
      wg_slot_id_gen_i <= _GEN_2;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_0_0 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (~cu_id_cancel & 2'h0 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_0_0 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_0_0 <= _GEN_24;
      end
    end else begin
      wg_slot_id_bitmap_0_0 <= _GEN_24;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_0_1 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (~cu_id_cancel & 2'h1 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_0_1 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_0_1 <= _GEN_25;
      end
    end else begin
      wg_slot_id_bitmap_0_1 <= _GEN_25;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_0_2 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (~cu_id_cancel & 2'h2 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_0_2 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_0_2 <= _GEN_26;
      end
    end else begin
      wg_slot_id_bitmap_0_2 <= _GEN_26;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_0_3 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (~cu_id_cancel & 2'h3 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_0_3 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_0_3 <= _GEN_27;
      end
    end else begin
      wg_slot_id_bitmap_0_3 <= _GEN_27;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_1_0 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (cu_id_cancel & 2'h0 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_1_0 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_1_0 <= _GEN_28;
      end
    end else begin
      wg_slot_id_bitmap_1_0 <= _GEN_28;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_1_1 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (cu_id_cancel & 2'h1 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_1_1 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_1_1 <= _GEN_29;
      end
    end else begin
      wg_slot_id_bitmap_1_1 <= _GEN_29;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_1_2 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (cu_id_cancel & 2'h2 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_1_2 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_1_2 <= _GEN_30;
      end
    end else begin
      wg_slot_id_bitmap_1_2 <= _GEN_30;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 20:36]
      wg_slot_id_bitmap_1_3 <= 1'h0; // @[wg_slot_id_convert_opt.scala 20:36]
    end else if (cancel_valid) begin // @[wg_slot_id_convert_opt.scala 80:23]
      if (cu_id_cancel & 2'h3 == wg_slot_id_find_i) begin // @[wg_slot_id_convert_opt.scala 81:60]
        wg_slot_id_bitmap_1_3 <= 1'h0; // @[wg_slot_id_convert_opt.scala 81:60]
      end else begin
        wg_slot_id_bitmap_1_3 <= _GEN_31;
      end
    end else begin
      wg_slot_id_bitmap_1_3 <= _GEN_31;
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_0_1 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (_GEN_72 & _GEN_76) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_0_1 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_0_2 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (_GEN_72 & _GEN_79) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_0_2 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_0_3 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (_GEN_72 & _GEN_82) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_0_3 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_1_0 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (io_cu_id & _GEN_73) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_1_0 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_1_1 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (io_cu_id & _GEN_76) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_1_1 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_1_2 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (io_cu_id & _GEN_79) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_1_2 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 52:42]
      wg_slot_id_find_ram_cam_1_3 <= 5'h0; // @[wg_slot_id_convert_opt.scala 52:42]
    end else if (_T_4) begin // @[wg_slot_id_convert_opt.scala 70:45]
      if (io_cu_id & _GEN_82) begin // @[wg_slot_id_convert_opt.scala 71:58]
        wg_slot_id_find_ram_cam_1_3 <= io_wg_id; // @[wg_slot_id_convert_opt.scala 71:58]
      end
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 75:31]
      cu_id_cancel <= 1'h0; // @[wg_slot_id_convert_opt.scala 75:31]
    end else begin
      cu_id_cancel <= io_cu_id; // @[wg_slot_id_convert_opt.scala 77:18]
    end
    if (reset) begin // @[wg_slot_id_convert_opt.scala 76:31]
      cancel_valid <= 1'h0; // @[wg_slot_id_convert_opt.scala 76:31]
    end else begin
      cancel_valid <= io_find_and_cancel; // @[wg_slot_id_convert_opt.scala 78:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wg_slot_id_find_i = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wg_slot_id_gen_i = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  wg_slot_id_bitmap_0_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wg_slot_id_bitmap_0_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wg_slot_id_bitmap_0_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wg_slot_id_bitmap_0_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  wg_slot_id_bitmap_1_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wg_slot_id_bitmap_1_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wg_slot_id_bitmap_1_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  wg_slot_id_bitmap_1_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_0_1 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_0_2 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_0_3 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_1_0 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_1_1 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_1_2 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  wg_slot_id_find_ram_cam_1_3 = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  cu_id_cancel = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  cancel_valid = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module throttling_engine(
  input        clock,
  input        reset,
  input        io_cu_id,
  input        io_alloc_en,
  input        io_dealloc_en,
  output [2:0] io_wg_count_available
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] actual_wg_count_array_0; // @[throttling_engine.scala 17:40]
  reg [2:0] actual_wg_count_array_1; // @[throttling_engine.scala 17:40]
  reg  cu_id_i; // @[throttling_engine.scala 26:26]
  reg  alloc_en_i; // @[throttling_engine.scala 27:29]
  reg  dealloc_en_i; // @[throttling_engine.scala 28:31]
  reg [2:0] wg_count_available_i; // @[throttling_engine.scala 34:39]
  wire [2:0] _GEN_10 = cu_id_i ? actual_wg_count_array_1 : actual_wg_count_array_0; // @[throttling_engine.scala 36:{38,38}]
  wire [2:0] _wg_count_available_i_T_1 = 3'h4 - _GEN_10; // @[throttling_engine.scala 37:61]
  wire [2:0] _actual_wg_count_array_T_1 = _GEN_10 + 3'h1; // @[throttling_engine.scala 43:74]
  wire [2:0] _GEN_12 = ~cu_id_i ? _actual_wg_count_array_T_1 : actual_wg_count_array_0; // @[throttling_engine.scala 17:40 43:{40,40}]
  wire [2:0] _GEN_13 = cu_id_i ? _actual_wg_count_array_T_1 : actual_wg_count_array_1; // @[throttling_engine.scala 17:40 43:{40,40}]
  wire [2:0] _GEN_14 = alloc_en_i ? _GEN_12 : actual_wg_count_array_0; // @[throttling_engine.scala 42:21 17:40]
  wire [2:0] _GEN_15 = alloc_en_i ? _GEN_13 : actual_wg_count_array_1; // @[throttling_engine.scala 42:21 17:40]
  wire [2:0] _actual_wg_count_array_T_3 = _GEN_10 - 3'h1; // @[throttling_engine.scala 46:74]
  assign io_wg_count_available = wg_count_available_i; // @[throttling_engine.scala 35:27]
  always @(posedge clock) begin
    if (reset) begin // @[throttling_engine.scala 17:40]
      actual_wg_count_array_0 <= 3'h0; // @[throttling_engine.scala 17:40]
    end else if (dealloc_en_i) begin // @[throttling_engine.scala 45:23]
      if (~cu_id_i) begin // @[throttling_engine.scala 46:40]
        actual_wg_count_array_0 <= _actual_wg_count_array_T_3; // @[throttling_engine.scala 46:40]
      end else begin
        actual_wg_count_array_0 <= _GEN_14;
      end
    end else begin
      actual_wg_count_array_0 <= _GEN_14;
    end
    if (reset) begin // @[throttling_engine.scala 17:40]
      actual_wg_count_array_1 <= 3'h0; // @[throttling_engine.scala 17:40]
    end else if (dealloc_en_i) begin // @[throttling_engine.scala 45:23]
      if (cu_id_i) begin // @[throttling_engine.scala 46:40]
        actual_wg_count_array_1 <= _actual_wg_count_array_T_3; // @[throttling_engine.scala 46:40]
      end else begin
        actual_wg_count_array_1 <= _GEN_15;
      end
    end else begin
      actual_wg_count_array_1 <= _GEN_15;
    end
    if (reset) begin // @[throttling_engine.scala 26:26]
      cu_id_i <= 1'h0; // @[throttling_engine.scala 26:26]
    end else if (io_alloc_en | io_dealloc_en) begin // @[throttling_engine.scala 31:39]
      cu_id_i <= io_cu_id; // @[throttling_engine.scala 32:17]
    end
    if (reset) begin // @[throttling_engine.scala 27:29]
      alloc_en_i <= 1'h0; // @[throttling_engine.scala 27:29]
    end else begin
      alloc_en_i <= io_alloc_en; // @[throttling_engine.scala 29:16]
    end
    if (reset) begin // @[throttling_engine.scala 28:31]
      dealloc_en_i <= 1'h0; // @[throttling_engine.scala 28:31]
    end else begin
      dealloc_en_i <= io_dealloc_en; // @[throttling_engine.scala 30:18]
    end
    if (reset) begin // @[throttling_engine.scala 34:39]
      wg_count_available_i <= 3'h0; // @[throttling_engine.scala 34:39]
    end else if (3'h4 > _GEN_10) begin // @[throttling_engine.scala 36:71]
      wg_count_available_i <= _wg_count_available_i_T_1; // @[throttling_engine.scala 37:30]
    end else begin
      wg_count_available_i <= 3'h0; // @[throttling_engine.scala 40:30]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  actual_wg_count_array_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  actual_wg_count_array_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  cu_id_i = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alloc_en_i = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dealloc_en_i = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wg_count_available_i = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module resource_table_group(
  input         clock,
  input         reset,
  input         io_alloc_en,
  input         io_dealloc_en,
  input  [4:0]  io_wg_id,
  input         io_sub_cu_id,
  output        io_res_tbl_done,
  output [12:0] io_lds_start,
  output [12:0] io_lds_size,
  output [12:0] io_vgpr_start,
  output [12:0] io_vgpr_size,
  output [12:0] io_sgpr_start,
  output [12:0] io_sgpr_size,
  output [2:0]  io_wf_count,
  output [2:0]  io_wg_count,
  input  [12:0] io_lds_start_in,
  input  [12:0] io_lds_size_in,
  input  [12:0] io_vgpr_start_in,
  input  [12:0] io_vgpr_size_in,
  input  [12:0] io_sgpr_start_in,
  input  [12:0] io_sgpr_size_in,
  input  [2:0]  io_wf_count_in,
  input         io_done_cancelled
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  lds_res_tbl_clock; // @[resource_table_group.scala 29:29]
  wire  lds_res_tbl_reset; // @[resource_table_group.scala 29:29]
  wire  lds_res_tbl_io_res_table_done_o; // @[resource_table_group.scala 29:29]
  wire [13:0] lds_res_tbl_io_cam_biggest_space_size; // @[resource_table_group.scala 29:29]
  wire [12:0] lds_res_tbl_io_cam_biggest_space_addr; // @[resource_table_group.scala 29:29]
  wire  lds_res_tbl_io_alloc_res_en; // @[resource_table_group.scala 29:29]
  wire  lds_res_tbl_io_dealloc_res_en; // @[resource_table_group.scala 29:29]
  wire  lds_res_tbl_io_alloc_cu_id; // @[resource_table_group.scala 29:29]
  wire  lds_res_tbl_io_dealloc_cu_id; // @[resource_table_group.scala 29:29]
  wire [1:0] lds_res_tbl_io_alloc_wg_slot_id; // @[resource_table_group.scala 29:29]
  wire [1:0] lds_res_tbl_io_dealloc_wg_slot_id; // @[resource_table_group.scala 29:29]
  wire [13:0] lds_res_tbl_io_alloc_res_size; // @[resource_table_group.scala 29:29]
  wire [12:0] lds_res_tbl_io_alloc_res_start; // @[resource_table_group.scala 29:29]
  wire  vgpr_res_tbl_clock; // @[resource_table_group.scala 30:30]
  wire  vgpr_res_tbl_reset; // @[resource_table_group.scala 30:30]
  wire  vgpr_res_tbl_io_res_table_done_o; // @[resource_table_group.scala 30:30]
  wire [13:0] vgpr_res_tbl_io_cam_biggest_space_size; // @[resource_table_group.scala 30:30]
  wire [12:0] vgpr_res_tbl_io_cam_biggest_space_addr; // @[resource_table_group.scala 30:30]
  wire  vgpr_res_tbl_io_alloc_res_en; // @[resource_table_group.scala 30:30]
  wire  vgpr_res_tbl_io_dealloc_res_en; // @[resource_table_group.scala 30:30]
  wire  vgpr_res_tbl_io_alloc_cu_id; // @[resource_table_group.scala 30:30]
  wire  vgpr_res_tbl_io_dealloc_cu_id; // @[resource_table_group.scala 30:30]
  wire [1:0] vgpr_res_tbl_io_alloc_wg_slot_id; // @[resource_table_group.scala 30:30]
  wire [1:0] vgpr_res_tbl_io_dealloc_wg_slot_id; // @[resource_table_group.scala 30:30]
  wire [13:0] vgpr_res_tbl_io_alloc_res_size; // @[resource_table_group.scala 30:30]
  wire [12:0] vgpr_res_tbl_io_alloc_res_start; // @[resource_table_group.scala 30:30]
  wire  sgpr_res_tbl_clock; // @[resource_table_group.scala 31:30]
  wire  sgpr_res_tbl_reset; // @[resource_table_group.scala 31:30]
  wire  sgpr_res_tbl_io_res_table_done_o; // @[resource_table_group.scala 31:30]
  wire [13:0] sgpr_res_tbl_io_cam_biggest_space_size; // @[resource_table_group.scala 31:30]
  wire [12:0] sgpr_res_tbl_io_cam_biggest_space_addr; // @[resource_table_group.scala 31:30]
  wire  sgpr_res_tbl_io_alloc_res_en; // @[resource_table_group.scala 31:30]
  wire  sgpr_res_tbl_io_dealloc_res_en; // @[resource_table_group.scala 31:30]
  wire  sgpr_res_tbl_io_alloc_cu_id; // @[resource_table_group.scala 31:30]
  wire  sgpr_res_tbl_io_dealloc_cu_id; // @[resource_table_group.scala 31:30]
  wire [1:0] sgpr_res_tbl_io_alloc_wg_slot_id; // @[resource_table_group.scala 31:30]
  wire [1:0] sgpr_res_tbl_io_dealloc_wg_slot_id; // @[resource_table_group.scala 31:30]
  wire [13:0] sgpr_res_tbl_io_alloc_res_size; // @[resource_table_group.scala 31:30]
  wire [12:0] sgpr_res_tbl_io_alloc_res_start; // @[resource_table_group.scala 31:30]
  wire  wf_res_tbl_clock; // @[resource_table_group.scala 32:28]
  wire  wf_res_tbl_reset; // @[resource_table_group.scala 32:28]
  wire [2:0] wf_res_tbl_io_wf_count_out; // @[resource_table_group.scala 32:28]
  wire  wf_res_tbl_io_cu_id; // @[resource_table_group.scala 32:28]
  wire  wf_res_tbl_io_alloc_en; // @[resource_table_group.scala 32:28]
  wire  wf_res_tbl_io_dealloc_en; // @[resource_table_group.scala 32:28]
  wire [2:0] wf_res_tbl_io_wf_count_in; // @[resource_table_group.scala 32:28]
  wire [1:0] wf_res_tbl_io_alloc_wg_slot_id; // @[resource_table_group.scala 32:28]
  wire [1:0] wf_res_tbl_io_dealloc_wg_slot_id; // @[resource_table_group.scala 32:28]
  wire  wf_slot_id_gen_clock; // @[resource_table_group.scala 33:32]
  wire  wf_slot_id_gen_reset; // @[resource_table_group.scala 33:32]
  wire [4:0] wf_slot_id_gen_io_wg_id; // @[resource_table_group.scala 33:32]
  wire  wf_slot_id_gen_io_cu_id; // @[resource_table_group.scala 33:32]
  wire [1:0] wf_slot_id_gen_io_wg_slot_id_gen; // @[resource_table_group.scala 33:32]
  wire [1:0] wf_slot_id_gen_io_wg_slot_id_find; // @[resource_table_group.scala 33:32]
  wire  wf_slot_id_gen_io_find_and_cancel; // @[resource_table_group.scala 33:32]
  wire  wf_slot_id_gen_io_generate; // @[resource_table_group.scala 33:32]
  wire  wg_throttling_clock; // @[resource_table_group.scala 34:31]
  wire  wg_throttling_reset; // @[resource_table_group.scala 34:31]
  wire  wg_throttling_io_cu_id; // @[resource_table_group.scala 34:31]
  wire  wg_throttling_io_alloc_en; // @[resource_table_group.scala 34:31]
  wire  wg_throttling_io_dealloc_en; // @[resource_table_group.scala 34:31]
  wire [2:0] wg_throttling_io_wg_count_available; // @[resource_table_group.scala 34:31]
  reg  alloc_en_1; // @[resource_table_group.scala 36:29]
  reg  dealloc_en_1; // @[resource_table_group.scala 38:31]
  reg  cu_id_1; // @[resource_table_group.scala 44:26]
  reg [12:0] lds_size1; // @[resource_table_group.scala 45:28]
  reg [12:0] vgpr_size1; // @[resource_table_group.scala 46:29]
  reg [12:0] sgpr_size1; // @[resource_table_group.scala 47:29]
  reg [2:0] wf_count1; // @[resource_table_group.scala 48:28]
  reg [12:0] lds_start1; // @[resource_table_group.scala 49:29]
  reg [12:0] vgpr_start1; // @[resource_table_group.scala 50:30]
  reg [12:0] sgpr_start1; // @[resource_table_group.scala 51:30]
  reg  lds_done_out; // @[resource_table_group.scala 52:31]
  reg  vgpr_done_out; // @[resource_table_group.scala 53:32]
  reg  sgpr_done_out; // @[resource_table_group.scala 54:32]
  wire  _GEN_7 = io_alloc_en | io_dealloc_en ? 1'h0 : lds_done_out; // @[resource_table_group.scala 57:39 65:22 52:31]
  wire  _GEN_8 = io_alloc_en | io_dealloc_en ? 1'h0 : vgpr_done_out; // @[resource_table_group.scala 57:39 66:23 53:32]
  wire  _GEN_9 = io_alloc_en | io_dealloc_en ? 1'h0 : sgpr_done_out; // @[resource_table_group.scala 57:39 67:23 54:32]
  reg [12:0] lds_size_out; // @[resource_table_group.scala 127:31]
  reg [12:0] vgpr_size_out; // @[resource_table_group.scala 128:32]
  reg [12:0] sgpr_size_out; // @[resource_table_group.scala 129:32]
  reg [12:0] lds_start_out; // @[resource_table_group.scala 130:32]
  reg [12:0] vgpr_start_out; // @[resource_table_group.scala 131:33]
  reg [12:0] sgpr_start_out; // @[resource_table_group.scala 132:33]
  wire  _GEN_12 = lds_res_tbl_io_res_table_done_o | _GEN_7; // @[resource_table_group.scala 133:42 134:22]
  wire [13:0] _GEN_13 = lds_res_tbl_io_res_table_done_o ? lds_res_tbl_io_cam_biggest_space_size : {{1'd0}, lds_size_out}
    ; // @[resource_table_group.scala 133:42 135:22 127:31]
  wire  _GEN_15 = vgpr_res_tbl_io_res_table_done_o | _GEN_8; // @[resource_table_group.scala 138:43 139:23]
  wire [13:0] _GEN_16 = vgpr_res_tbl_io_res_table_done_o ? vgpr_res_tbl_io_cam_biggest_space_size : {{1'd0},
    vgpr_size_out}; // @[resource_table_group.scala 138:43 140:23 128:32]
  wire  _GEN_18 = sgpr_res_tbl_io_res_table_done_o | _GEN_9; // @[resource_table_group.scala 143:43 144:23]
  wire [13:0] _GEN_19 = sgpr_res_tbl_io_res_table_done_o ? sgpr_res_tbl_io_cam_biggest_space_size : {{1'd0},
    sgpr_size_out}; // @[resource_table_group.scala 143:43 145:23 129:32]
  wire [13:0] _GEN_24 = reset ? 14'h0 : _GEN_13; // @[resource_table_group.scala 127:{31,31}]
  wire [13:0] _GEN_25 = reset ? 14'h0 : _GEN_16; // @[resource_table_group.scala 128:{32,32}]
  wire [13:0] _GEN_26 = reset ? 14'h0 : _GEN_19; // @[resource_table_group.scala 129:{32,32}]
  resource_table lds_res_tbl ( // @[resource_table_group.scala 29:29]
    .clock(lds_res_tbl_clock),
    .reset(lds_res_tbl_reset),
    .io_res_table_done_o(lds_res_tbl_io_res_table_done_o),
    .io_cam_biggest_space_size(lds_res_tbl_io_cam_biggest_space_size),
    .io_cam_biggest_space_addr(lds_res_tbl_io_cam_biggest_space_addr),
    .io_alloc_res_en(lds_res_tbl_io_alloc_res_en),
    .io_dealloc_res_en(lds_res_tbl_io_dealloc_res_en),
    .io_alloc_cu_id(lds_res_tbl_io_alloc_cu_id),
    .io_dealloc_cu_id(lds_res_tbl_io_dealloc_cu_id),
    .io_alloc_wg_slot_id(lds_res_tbl_io_alloc_wg_slot_id),
    .io_dealloc_wg_slot_id(lds_res_tbl_io_dealloc_wg_slot_id),
    .io_alloc_res_size(lds_res_tbl_io_alloc_res_size),
    .io_alloc_res_start(lds_res_tbl_io_alloc_res_start)
  );
  resource_table vgpr_res_tbl ( // @[resource_table_group.scala 30:30]
    .clock(vgpr_res_tbl_clock),
    .reset(vgpr_res_tbl_reset),
    .io_res_table_done_o(vgpr_res_tbl_io_res_table_done_o),
    .io_cam_biggest_space_size(vgpr_res_tbl_io_cam_biggest_space_size),
    .io_cam_biggest_space_addr(vgpr_res_tbl_io_cam_biggest_space_addr),
    .io_alloc_res_en(vgpr_res_tbl_io_alloc_res_en),
    .io_dealloc_res_en(vgpr_res_tbl_io_dealloc_res_en),
    .io_alloc_cu_id(vgpr_res_tbl_io_alloc_cu_id),
    .io_dealloc_cu_id(vgpr_res_tbl_io_dealloc_cu_id),
    .io_alloc_wg_slot_id(vgpr_res_tbl_io_alloc_wg_slot_id),
    .io_dealloc_wg_slot_id(vgpr_res_tbl_io_dealloc_wg_slot_id),
    .io_alloc_res_size(vgpr_res_tbl_io_alloc_res_size),
    .io_alloc_res_start(vgpr_res_tbl_io_alloc_res_start)
  );
  resource_table sgpr_res_tbl ( // @[resource_table_group.scala 31:30]
    .clock(sgpr_res_tbl_clock),
    .reset(sgpr_res_tbl_reset),
    .io_res_table_done_o(sgpr_res_tbl_io_res_table_done_o),
    .io_cam_biggest_space_size(sgpr_res_tbl_io_cam_biggest_space_size),
    .io_cam_biggest_space_addr(sgpr_res_tbl_io_cam_biggest_space_addr),
    .io_alloc_res_en(sgpr_res_tbl_io_alloc_res_en),
    .io_dealloc_res_en(sgpr_res_tbl_io_dealloc_res_en),
    .io_alloc_cu_id(sgpr_res_tbl_io_alloc_cu_id),
    .io_dealloc_cu_id(sgpr_res_tbl_io_dealloc_cu_id),
    .io_alloc_wg_slot_id(sgpr_res_tbl_io_alloc_wg_slot_id),
    .io_dealloc_wg_slot_id(sgpr_res_tbl_io_dealloc_wg_slot_id),
    .io_alloc_res_size(sgpr_res_tbl_io_alloc_res_size),
    .io_alloc_res_start(sgpr_res_tbl_io_alloc_res_start)
  );
  wg_resource_table_neo wf_res_tbl ( // @[resource_table_group.scala 32:28]
    .clock(wf_res_tbl_clock),
    .reset(wf_res_tbl_reset),
    .io_wf_count_out(wf_res_tbl_io_wf_count_out),
    .io_cu_id(wf_res_tbl_io_cu_id),
    .io_alloc_en(wf_res_tbl_io_alloc_en),
    .io_dealloc_en(wf_res_tbl_io_dealloc_en),
    .io_wf_count_in(wf_res_tbl_io_wf_count_in),
    .io_alloc_wg_slot_id(wf_res_tbl_io_alloc_wg_slot_id),
    .io_dealloc_wg_slot_id(wf_res_tbl_io_dealloc_wg_slot_id)
  );
  wg_slot_id_convert_opt wf_slot_id_gen ( // @[resource_table_group.scala 33:32]
    .clock(wf_slot_id_gen_clock),
    .reset(wf_slot_id_gen_reset),
    .io_wg_id(wf_slot_id_gen_io_wg_id),
    .io_cu_id(wf_slot_id_gen_io_cu_id),
    .io_wg_slot_id_gen(wf_slot_id_gen_io_wg_slot_id_gen),
    .io_wg_slot_id_find(wf_slot_id_gen_io_wg_slot_id_find),
    .io_find_and_cancel(wf_slot_id_gen_io_find_and_cancel),
    .io_generate(wf_slot_id_gen_io_generate)
  );
  throttling_engine wg_throttling ( // @[resource_table_group.scala 34:31]
    .clock(wg_throttling_clock),
    .reset(wg_throttling_reset),
    .io_cu_id(wg_throttling_io_cu_id),
    .io_alloc_en(wg_throttling_io_alloc_en),
    .io_dealloc_en(wg_throttling_io_dealloc_en),
    .io_wg_count_available(wg_throttling_io_wg_count_available)
  );
  assign io_res_tbl_done = lds_done_out & vgpr_done_out & sgpr_done_out; // @[resource_table_group.scala 56:54]
  assign io_lds_start = lds_start_out; // @[resource_table_group.scala 151:18]
  assign io_lds_size = lds_size_out; // @[resource_table_group.scala 148:17]
  assign io_vgpr_start = vgpr_start_out; // @[resource_table_group.scala 152:19]
  assign io_vgpr_size = vgpr_size_out; // @[resource_table_group.scala 149:18]
  assign io_sgpr_start = sgpr_start_out; // @[resource_table_group.scala 153:19]
  assign io_sgpr_size = sgpr_size_out; // @[resource_table_group.scala 150:18]
  assign io_wf_count = wf_res_tbl_io_wf_count_out; // @[resource_table_group.scala 125:17]
  assign io_wg_count = wg_throttling_io_wg_count_available; // @[resource_table_group.scala 126:17]
  assign lds_res_tbl_clock = clock;
  assign lds_res_tbl_reset = reset;
  assign lds_res_tbl_io_alloc_res_en = alloc_en_1; // @[resource_table_group.scala 77:33]
  assign lds_res_tbl_io_dealloc_res_en = dealloc_en_1; // @[resource_table_group.scala 78:35]
  assign lds_res_tbl_io_alloc_cu_id = cu_id_1; // @[resource_table_group.scala 79:32]
  assign lds_res_tbl_io_dealloc_cu_id = cu_id_1; // @[resource_table_group.scala 80:34]
  assign lds_res_tbl_io_alloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_gen; // @[resource_table_group.scala 81:37]
  assign lds_res_tbl_io_dealloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_find; // @[resource_table_group.scala 82:39]
  assign lds_res_tbl_io_alloc_res_size = {{1'd0}, lds_size1}; // @[resource_table_group.scala 83:35]
  assign lds_res_tbl_io_alloc_res_start = lds_start1; // @[resource_table_group.scala 84:36]
  assign vgpr_res_tbl_clock = clock;
  assign vgpr_res_tbl_reset = reset;
  assign vgpr_res_tbl_io_alloc_res_en = alloc_en_1; // @[resource_table_group.scala 86:34]
  assign vgpr_res_tbl_io_dealloc_res_en = dealloc_en_1; // @[resource_table_group.scala 87:36]
  assign vgpr_res_tbl_io_alloc_cu_id = cu_id_1; // @[resource_table_group.scala 88:33]
  assign vgpr_res_tbl_io_dealloc_cu_id = cu_id_1; // @[resource_table_group.scala 89:35]
  assign vgpr_res_tbl_io_alloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_gen; // @[resource_table_group.scala 90:38]
  assign vgpr_res_tbl_io_dealloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_find; // @[resource_table_group.scala 91:40]
  assign vgpr_res_tbl_io_alloc_res_size = {{1'd0}, vgpr_size1}; // @[resource_table_group.scala 92:36]
  assign vgpr_res_tbl_io_alloc_res_start = vgpr_start1; // @[resource_table_group.scala 93:37]
  assign sgpr_res_tbl_clock = clock;
  assign sgpr_res_tbl_reset = reset;
  assign sgpr_res_tbl_io_alloc_res_en = alloc_en_1; // @[resource_table_group.scala 95:34]
  assign sgpr_res_tbl_io_dealloc_res_en = dealloc_en_1; // @[resource_table_group.scala 96:36]
  assign sgpr_res_tbl_io_alloc_cu_id = cu_id_1; // @[resource_table_group.scala 97:33]
  assign sgpr_res_tbl_io_dealloc_cu_id = cu_id_1; // @[resource_table_group.scala 98:35]
  assign sgpr_res_tbl_io_alloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_gen; // @[resource_table_group.scala 99:38]
  assign sgpr_res_tbl_io_dealloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_find; // @[resource_table_group.scala 100:40]
  assign sgpr_res_tbl_io_alloc_res_size = {{1'd0}, sgpr_size1}; // @[resource_table_group.scala 101:36]
  assign sgpr_res_tbl_io_alloc_res_start = sgpr_start1; // @[resource_table_group.scala 102:37]
  assign wf_res_tbl_clock = clock;
  assign wf_res_tbl_reset = reset;
  assign wf_res_tbl_io_cu_id = cu_id_1; // @[resource_table_group.scala 104:25]
  assign wf_res_tbl_io_alloc_en = alloc_en_1; // @[resource_table_group.scala 105:28]
  assign wf_res_tbl_io_dealloc_en = dealloc_en_1; // @[resource_table_group.scala 106:30]
  assign wf_res_tbl_io_wf_count_in = wf_count1; // @[resource_table_group.scala 107:31]
  assign wf_res_tbl_io_alloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_gen; // @[resource_table_group.scala 108:36]
  assign wf_res_tbl_io_dealloc_wg_slot_id = wf_slot_id_gen_io_wg_slot_id_find; // @[resource_table_group.scala 109:38]
  assign wf_slot_id_gen_clock = clock;
  assign wf_slot_id_gen_reset = reset;
  assign wf_slot_id_gen_io_wg_id = io_wg_id; // @[resource_table_group.scala 40:29]
  assign wf_slot_id_gen_io_cu_id = io_sub_cu_id; // @[resource_table_group.scala 41:29]
  assign wf_slot_id_gen_io_find_and_cancel = io_dealloc_en; // @[resource_table_group.scala 43:39]
  assign wf_slot_id_gen_io_generate = io_alloc_en; // @[resource_table_group.scala 42:32]
  assign wg_throttling_clock = clock;
  assign wg_throttling_reset = reset;
  assign wg_throttling_io_cu_id = cu_id_1; // @[resource_table_group.scala 111:28]
  assign wg_throttling_io_alloc_en = alloc_en_1; // @[resource_table_group.scala 112:31]
  assign wg_throttling_io_dealloc_en = dealloc_en_1; // @[resource_table_group.scala 113:33]
  always @(posedge clock) begin
    if (reset) begin // @[resource_table_group.scala 36:29]
      alloc_en_1 <= 1'h0; // @[resource_table_group.scala 36:29]
    end else begin
      alloc_en_1 <= io_alloc_en; // @[resource_table_group.scala 37:16]
    end
    if (reset) begin // @[resource_table_group.scala 38:31]
      dealloc_en_1 <= 1'h0; // @[resource_table_group.scala 38:31]
    end else begin
      dealloc_en_1 <= io_dealloc_en; // @[resource_table_group.scala 39:18]
    end
    if (reset) begin // @[resource_table_group.scala 44:26]
      cu_id_1 <= 1'h0; // @[resource_table_group.scala 44:26]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      cu_id_1 <= io_sub_cu_id; // @[resource_table_group.scala 58:17]
    end
    if (reset) begin // @[resource_table_group.scala 45:28]
      lds_size1 <= 13'h0; // @[resource_table_group.scala 45:28]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      lds_size1 <= io_lds_size_in; // @[resource_table_group.scala 59:19]
    end
    if (reset) begin // @[resource_table_group.scala 46:29]
      vgpr_size1 <= 13'h0; // @[resource_table_group.scala 46:29]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      vgpr_size1 <= io_vgpr_size_in; // @[resource_table_group.scala 60:20]
    end
    if (reset) begin // @[resource_table_group.scala 47:29]
      sgpr_size1 <= 13'h0; // @[resource_table_group.scala 47:29]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      sgpr_size1 <= io_sgpr_size_in; // @[resource_table_group.scala 61:20]
    end
    if (reset) begin // @[resource_table_group.scala 48:28]
      wf_count1 <= 3'h0; // @[resource_table_group.scala 48:28]
    end else if (io_alloc_en) begin // @[resource_table_group.scala 69:22]
      wf_count1 <= io_wf_count_in; // @[resource_table_group.scala 70:19]
    end else if (io_dealloc_en) begin // @[resource_table_group.scala 73:29]
      wf_count1 <= 3'h0; // @[resource_table_group.scala 74:19]
    end
    if (reset) begin // @[resource_table_group.scala 49:29]
      lds_start1 <= 13'h0; // @[resource_table_group.scala 49:29]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      lds_start1 <= io_lds_start_in; // @[resource_table_group.scala 62:20]
    end
    if (reset) begin // @[resource_table_group.scala 50:30]
      vgpr_start1 <= 13'h0; // @[resource_table_group.scala 50:30]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      vgpr_start1 <= io_vgpr_start_in; // @[resource_table_group.scala 63:21]
    end
    if (reset) begin // @[resource_table_group.scala 51:30]
      sgpr_start1 <= 13'h0; // @[resource_table_group.scala 51:30]
    end else if (io_alloc_en | io_dealloc_en) begin // @[resource_table_group.scala 57:39]
      sgpr_start1 <= io_sgpr_start_in; // @[resource_table_group.scala 64:21]
    end
    if (reset) begin // @[resource_table_group.scala 52:31]
      lds_done_out <= 1'h0; // @[resource_table_group.scala 52:31]
    end else if (io_done_cancelled) begin // @[resource_table_group.scala 154:28]
      lds_done_out <= 1'h0; // @[resource_table_group.scala 156:22]
    end else begin
      lds_done_out <= _GEN_12;
    end
    if (reset) begin // @[resource_table_group.scala 53:32]
      vgpr_done_out <= 1'h0; // @[resource_table_group.scala 53:32]
    end else if (io_done_cancelled) begin // @[resource_table_group.scala 154:28]
      vgpr_done_out <= 1'h0; // @[resource_table_group.scala 157:23]
    end else begin
      vgpr_done_out <= _GEN_15;
    end
    if (reset) begin // @[resource_table_group.scala 54:32]
      sgpr_done_out <= 1'h0; // @[resource_table_group.scala 54:32]
    end else if (io_done_cancelled) begin // @[resource_table_group.scala 154:28]
      sgpr_done_out <= 1'h0; // @[resource_table_group.scala 158:23]
    end else begin
      sgpr_done_out <= _GEN_18;
    end
    lds_size_out <= _GEN_24[12:0]; // @[resource_table_group.scala 127:{31,31}]
    vgpr_size_out <= _GEN_25[12:0]; // @[resource_table_group.scala 128:{32,32}]
    sgpr_size_out <= _GEN_26[12:0]; // @[resource_table_group.scala 129:{32,32}]
    if (reset) begin // @[resource_table_group.scala 130:32]
      lds_start_out <= 13'h0; // @[resource_table_group.scala 130:32]
    end else if (lds_res_tbl_io_res_table_done_o) begin // @[resource_table_group.scala 133:42]
      lds_start_out <= lds_res_tbl_io_cam_biggest_space_addr; // @[resource_table_group.scala 136:23]
    end
    if (reset) begin // @[resource_table_group.scala 131:33]
      vgpr_start_out <= 13'h0; // @[resource_table_group.scala 131:33]
    end else if (vgpr_res_tbl_io_res_table_done_o) begin // @[resource_table_group.scala 138:43]
      vgpr_start_out <= vgpr_res_tbl_io_cam_biggest_space_addr; // @[resource_table_group.scala 141:24]
    end
    if (reset) begin // @[resource_table_group.scala 132:33]
      sgpr_start_out <= 13'h0; // @[resource_table_group.scala 132:33]
    end else if (sgpr_res_tbl_io_res_table_done_o) begin // @[resource_table_group.scala 143:43]
      sgpr_start_out <= sgpr_res_tbl_io_cam_biggest_space_addr; // @[resource_table_group.scala 146:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  alloc_en_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dealloc_en_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cu_id_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lds_size1 = _RAND_3[12:0];
  _RAND_4 = {1{`RANDOM}};
  vgpr_size1 = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  sgpr_size1 = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  wf_count1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  lds_start1 = _RAND_7[12:0];
  _RAND_8 = {1{`RANDOM}};
  vgpr_start1 = _RAND_8[12:0];
  _RAND_9 = {1{`RANDOM}};
  sgpr_start1 = _RAND_9[12:0];
  _RAND_10 = {1{`RANDOM}};
  lds_done_out = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vgpr_done_out = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  sgpr_done_out = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lds_size_out = _RAND_13[12:0];
  _RAND_14 = {1{`RANDOM}};
  vgpr_size_out = _RAND_14[12:0];
  _RAND_15 = {1{`RANDOM}};
  sgpr_size_out = _RAND_15[12:0];
  _RAND_16 = {1{`RANDOM}};
  lds_start_out = _RAND_16[12:0];
  _RAND_17 = {1{`RANDOM}};
  vgpr_start_out = _RAND_17[12:0];
  _RAND_18 = {1{`RANDOM}};
  sgpr_start_out = _RAND_18[12:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top_resource_table(
  input         clock,
  input         reset,
  output        io_grt_cam_up_valid,
  output [2:0]  io_grt_cam_up_wf_count,
  output [1:0]  io_grt_cam_up_cu_id,
  output [11:0] io_grt_cam_up_vgpr_strt,
  output [12:0] io_grt_cam_up_vgpr_size,
  output [11:0] io_grt_cam_up_sgpr_strt,
  output [12:0] io_grt_cam_up_sgpr_size,
  output [11:0] io_grt_cam_up_lds_strt,
  output [12:0] io_grt_cam_up_lds_size,
  output [2:0]  io_grt_cam_up_wg_count,
  output        io_grt_wg_alloc_done,
  output [1:0]  io_grt_wg_alloc_cu_id,
  output        io_grt_wg_dealloc_done,
  output [1:0]  io_grt_wg_dealloc_cu_id,
  input  [1:0]  io_gpu_interface_cu_id,
  input  [4:0]  io_gpu_interface_dealloc_wg_id,
  input         io_dis_controller_wg_alloc_valid,
  input         io_dis_controller_wg_dealloc_valid,
  input  [4:0]  io_allocator_wg_id_out,
  input  [2:0]  io_allocator_wf_count,
  input  [1:0]  io_allocator_cu_id_out,
  input  [11:0] io_allocator_vgpr_start_out,
  input  [12:0] io_allocator_vgpr_size_out,
  input  [11:0] io_allocator_sgpr_start_out,
  input  [12:0] io_allocator_sgpr_size_out,
  input  [11:0] io_allocator_lds_start_out,
  input  [12:0] io_allocator_lds_size_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  rt_group_clock; // @[top_resource_table.scala 54:30]
  wire  rt_group_reset; // @[top_resource_table.scala 54:30]
  wire  rt_group_io_alloc_en; // @[top_resource_table.scala 54:30]
  wire  rt_group_io_dealloc_en; // @[top_resource_table.scala 54:30]
  wire [4:0] rt_group_io_wg_id; // @[top_resource_table.scala 54:30]
  wire  rt_group_io_sub_cu_id; // @[top_resource_table.scala 54:30]
  wire  rt_group_io_res_tbl_done; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_lds_start; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_lds_size; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_vgpr_start; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_vgpr_size; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_sgpr_start; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_sgpr_size; // @[top_resource_table.scala 54:30]
  wire [2:0] rt_group_io_wf_count; // @[top_resource_table.scala 54:30]
  wire [2:0] rt_group_io_wg_count; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_lds_start_in; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_lds_size_in; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_vgpr_start_in; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_vgpr_size_in; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_sgpr_start_in; // @[top_resource_table.scala 54:30]
  wire [12:0] rt_group_io_sgpr_size_in; // @[top_resource_table.scala 54:30]
  wire [2:0] rt_group_io_wf_count_in; // @[top_resource_table.scala 54:30]
  wire  rt_group_io_done_cancelled; // @[top_resource_table.scala 54:30]
  reg  done_array_0; // @[top_resource_table.scala 38:29]
  reg [2:0] wf_count_array_0; // @[top_resource_table.scala 39:33]
  reg [2:0] wg_count_array_0; // @[top_resource_table.scala 40:33]
  reg [12:0] vgpr_start_array_0; // @[top_resource_table.scala 41:35]
  reg [12:0] vgpr_size_array_0; // @[top_resource_table.scala 42:34]
  reg [12:0] sgpr_start_array_0; // @[top_resource_table.scala 43:35]
  reg [12:0] sgpr_size_array_0; // @[top_resource_table.scala 44:34]
  reg [12:0] lds_start_array_0; // @[top_resource_table.scala 45:34]
  reg [12:0] lds_size_array_0; // @[top_resource_table.scala 46:33]
  reg [1:0] cu_id_array_0; // @[top_resource_table.scala 48:30]
  reg  serviced_array_0; // @[top_resource_table.scala 49:33]
  reg  is_alloc_array_0; // @[top_resource_table.scala 50:33]
  reg  done_cancelled_array_0; // @[top_resource_table.scala 51:39]
  reg  command_serviced_array_cancelled_0; // @[top_resource_table.scala 52:51]
  wire  _GEN_5 = io_dis_controller_wg_alloc_valid & ~io_allocator_cu_id_out[1] | command_serviced_array_cancelled_0; // @[top_resource_table.scala 71:134 75:49 52:51]
  wire  _GEN_6 = io_dis_controller_wg_alloc_valid & ~io_allocator_cu_id_out[1] ? 1'h0 : done_cancelled_array_0; // @[top_resource_table.scala 71:134 76:37 51:39]
  wire  _GEN_7 = io_dis_controller_wg_alloc_valid & ~io_allocator_cu_id_out[1] | is_alloc_array_0; // @[top_resource_table.scala 71:134 77:31 50:33]
  wire  _GEN_11 = io_dis_controller_wg_dealloc_valid & ~io_gpu_interface_cu_id[1] | _GEN_5; // @[top_resource_table.scala 82:136 86:49]
  wire  _GEN_12 = io_dis_controller_wg_dealloc_valid & ~io_gpu_interface_cu_id[1] ? 1'h0 : _GEN_6; // @[top_resource_table.scala 82:136 87:37]
  wire  _GEN_14 = command_serviced_array_cancelled_0 ? 1'h0 : serviced_array_0; // @[top_resource_table.scala 102:50 103:31 49:33]
  wire  serviced_id_valid = done_array_0 & ~serviced_array_0; // @[top_resource_table.scala 114:28]
  reg  grt_cam_up_valid_i; // @[top_resource_table.scala 134:37]
  reg  grt_wg_alloc_done; // @[top_resource_table.scala 135:36]
  reg  grt_wg_dealloc_done; // @[top_resource_table.scala 136:38]
  wire  _GEN_19 = is_alloc_array_0 ? 1'h0 : 1'h1; // @[top_resource_table.scala 142:42 144:33 147:33]
  wire  _GEN_20 = serviced_id_valid | _GEN_14; // @[top_resource_table.scala 137:28 138:37]
  wire  _GEN_22 = serviced_id_valid | _GEN_12; // @[top_resource_table.scala 137:28 140:43]
  wire  _GEN_23 = serviced_id_valid & is_alloc_array_0; // @[top_resource_table.scala 137:28 153:27]
  wire  _GEN_24 = serviced_id_valid & _GEN_19; // @[top_resource_table.scala 137:28 154:29]
  resource_table_group rt_group ( // @[top_resource_table.scala 54:30]
    .clock(rt_group_clock),
    .reset(rt_group_reset),
    .io_alloc_en(rt_group_io_alloc_en),
    .io_dealloc_en(rt_group_io_dealloc_en),
    .io_wg_id(rt_group_io_wg_id),
    .io_sub_cu_id(rt_group_io_sub_cu_id),
    .io_res_tbl_done(rt_group_io_res_tbl_done),
    .io_lds_start(rt_group_io_lds_start),
    .io_lds_size(rt_group_io_lds_size),
    .io_vgpr_start(rt_group_io_vgpr_start),
    .io_vgpr_size(rt_group_io_vgpr_size),
    .io_sgpr_start(rt_group_io_sgpr_start),
    .io_sgpr_size(rt_group_io_sgpr_size),
    .io_wf_count(rt_group_io_wf_count),
    .io_wg_count(rt_group_io_wg_count),
    .io_lds_start_in(rt_group_io_lds_start_in),
    .io_lds_size_in(rt_group_io_lds_size_in),
    .io_vgpr_start_in(rt_group_io_vgpr_start_in),
    .io_vgpr_size_in(rt_group_io_vgpr_size_in),
    .io_sgpr_start_in(rt_group_io_sgpr_start_in),
    .io_sgpr_size_in(rt_group_io_sgpr_size_in),
    .io_wf_count_in(rt_group_io_wf_count_in),
    .io_done_cancelled(rt_group_io_done_cancelled)
  );
  assign io_grt_cam_up_valid = grt_cam_up_valid_i; // @[top_resource_table.scala 156:25]
  assign io_grt_cam_up_wf_count = wf_count_array_0; // @[top_resource_table.scala 127:28]
  assign io_grt_cam_up_cu_id = cu_id_array_0; // @[top_resource_table.scala 129:25]
  assign io_grt_cam_up_vgpr_strt = vgpr_start_array_0[11:0]; // @[top_resource_table.scala 121:29]
  assign io_grt_cam_up_vgpr_size = vgpr_size_array_0; // @[top_resource_table.scala 122:29]
  assign io_grt_cam_up_sgpr_strt = sgpr_start_array_0[11:0]; // @[top_resource_table.scala 123:29]
  assign io_grt_cam_up_sgpr_size = sgpr_size_array_0; // @[top_resource_table.scala 124:29]
  assign io_grt_cam_up_lds_strt = lds_start_array_0[11:0]; // @[top_resource_table.scala 125:28]
  assign io_grt_cam_up_lds_size = lds_size_array_0; // @[top_resource_table.scala 126:28]
  assign io_grt_cam_up_wg_count = wg_count_array_0; // @[top_resource_table.scala 128:28]
  assign io_grt_wg_alloc_done = grt_wg_alloc_done; // @[top_resource_table.scala 157:26]
  assign io_grt_wg_alloc_cu_id = cu_id_array_0; // @[top_resource_table.scala 130:27]
  assign io_grt_wg_dealloc_done = grt_wg_dealloc_done; // @[top_resource_table.scala 158:28]
  assign io_grt_wg_dealloc_cu_id = cu_id_array_0; // @[top_resource_table.scala 132:29]
  assign rt_group_clock = clock;
  assign rt_group_reset = reset;
  assign rt_group_io_alloc_en = io_dis_controller_wg_alloc_valid & ~io_allocator_cu_id_out[1]; // @[top_resource_table.scala 71:47]
  assign rt_group_io_dealloc_en = io_dis_controller_wg_dealloc_valid & ~io_gpu_interface_cu_id[1]; // @[top_resource_table.scala 82:49]
  assign rt_group_io_wg_id = io_dis_controller_wg_alloc_valid ? io_allocator_wg_id_out : io_gpu_interface_dealloc_wg_id; // @[top_resource_table.scala 63:47 64:31 68:31]
  assign rt_group_io_sub_cu_id = io_dis_controller_wg_alloc_valid ? io_allocator_cu_id_out[0] : io_gpu_interface_cu_id[0
    ]; // @[top_resource_table.scala 63:47 65:35 69:35]
  assign rt_group_io_lds_start_in = {1'h0,io_allocator_lds_start_out}; // @[Cat.scala 31:58]
  assign rt_group_io_lds_size_in = io_allocator_lds_size_out; // @[top_resource_table.scala 56:33]
  assign rt_group_io_vgpr_start_in = {1'h0,io_allocator_vgpr_start_out}; // @[Cat.scala 31:58]
  assign rt_group_io_vgpr_size_in = io_allocator_vgpr_size_out; // @[top_resource_table.scala 58:34]
  assign rt_group_io_sgpr_start_in = {1'h0,io_allocator_sgpr_start_out}; // @[Cat.scala 31:58]
  assign rt_group_io_sgpr_size_in = io_allocator_sgpr_size_out; // @[top_resource_table.scala 60:34]
  assign rt_group_io_wf_count_in = io_allocator_wf_count; // @[top_resource_table.scala 61:33]
  assign rt_group_io_done_cancelled = done_cancelled_array_0; // @[top_resource_table.scala 62:36]
  always @(posedge clock) begin
    if (reset) begin // @[top_resource_table.scala 38:29]
      done_array_0 <= 1'h0; // @[top_resource_table.scala 38:29]
    end else begin
      done_array_0 <= rt_group_io_res_tbl_done; // @[top_resource_table.scala 93:23]
    end
    if (reset) begin // @[top_resource_table.scala 39:33]
      wf_count_array_0 <= 3'h0; // @[top_resource_table.scala 39:33]
    end else begin
      wf_count_array_0 <= rt_group_io_wf_count; // @[top_resource_table.scala 94:27]
    end
    if (reset) begin // @[top_resource_table.scala 40:33]
      wg_count_array_0 <= 3'h0; // @[top_resource_table.scala 40:33]
    end else begin
      wg_count_array_0 <= rt_group_io_wg_count; // @[top_resource_table.scala 95:27]
    end
    if (reset) begin // @[top_resource_table.scala 41:35]
      vgpr_start_array_0 <= 13'h0; // @[top_resource_table.scala 41:35]
    end else begin
      vgpr_start_array_0 <= rt_group_io_vgpr_start; // @[top_resource_table.scala 96:29]
    end
    if (reset) begin // @[top_resource_table.scala 42:34]
      vgpr_size_array_0 <= 13'h0; // @[top_resource_table.scala 42:34]
    end else begin
      vgpr_size_array_0 <= rt_group_io_vgpr_size; // @[top_resource_table.scala 97:28]
    end
    if (reset) begin // @[top_resource_table.scala 43:35]
      sgpr_start_array_0 <= 13'h0; // @[top_resource_table.scala 43:35]
    end else begin
      sgpr_start_array_0 <= rt_group_io_sgpr_start; // @[top_resource_table.scala 98:29]
    end
    if (reset) begin // @[top_resource_table.scala 44:34]
      sgpr_size_array_0 <= 13'h0; // @[top_resource_table.scala 44:34]
    end else begin
      sgpr_size_array_0 <= rt_group_io_sgpr_size; // @[top_resource_table.scala 99:28]
    end
    if (reset) begin // @[top_resource_table.scala 45:34]
      lds_start_array_0 <= 13'h0; // @[top_resource_table.scala 45:34]
    end else begin
      lds_start_array_0 <= rt_group_io_lds_start; // @[top_resource_table.scala 100:28]
    end
    if (reset) begin // @[top_resource_table.scala 46:33]
      lds_size_array_0 <= 13'h0; // @[top_resource_table.scala 46:33]
    end else begin
      lds_size_array_0 <= rt_group_io_lds_size; // @[top_resource_table.scala 101:27]
    end
    if (reset) begin // @[top_resource_table.scala 48:30]
      cu_id_array_0 <= 2'h0; // @[top_resource_table.scala 48:30]
    end else if (io_dis_controller_wg_dealloc_valid & ~io_gpu_interface_cu_id[1]) begin // @[top_resource_table.scala 82:136]
      cu_id_array_0 <= io_gpu_interface_cu_id; // @[top_resource_table.scala 85:28]
    end else if (io_dis_controller_wg_alloc_valid & ~io_allocator_cu_id_out[1]) begin // @[top_resource_table.scala 71:134]
      cu_id_array_0 <= io_allocator_cu_id_out; // @[top_resource_table.scala 74:28]
    end
    if (reset) begin // @[top_resource_table.scala 49:33]
      serviced_array_0 <= 1'h0; // @[top_resource_table.scala 49:33]
    end else begin
      serviced_array_0 <= _GEN_20;
    end
    if (reset) begin // @[top_resource_table.scala 50:33]
      is_alloc_array_0 <= 1'h0; // @[top_resource_table.scala 50:33]
    end else if (io_dis_controller_wg_dealloc_valid & ~io_gpu_interface_cu_id[1]) begin // @[top_resource_table.scala 82:136]
      is_alloc_array_0 <= 1'h0; // @[top_resource_table.scala 88:31]
    end else begin
      is_alloc_array_0 <= _GEN_7;
    end
    if (reset) begin // @[top_resource_table.scala 51:39]
      done_cancelled_array_0 <= 1'h0; // @[top_resource_table.scala 51:39]
    end else begin
      done_cancelled_array_0 <= _GEN_22;
    end
    if (reset) begin // @[top_resource_table.scala 52:51]
      command_serviced_array_cancelled_0 <= 1'h0; // @[top_resource_table.scala 52:51]
    end else if (command_serviced_array_cancelled_0) begin // @[top_resource_table.scala 102:50]
      command_serviced_array_cancelled_0 <= 1'h0; // @[top_resource_table.scala 104:49]
    end else begin
      command_serviced_array_cancelled_0 <= _GEN_11;
    end
    if (reset) begin // @[top_resource_table.scala 134:37]
      grt_cam_up_valid_i <= 1'h0; // @[top_resource_table.scala 134:37]
    end else begin
      grt_cam_up_valid_i <= serviced_id_valid;
    end
    if (reset) begin // @[top_resource_table.scala 135:36]
      grt_wg_alloc_done <= 1'h0; // @[top_resource_table.scala 135:36]
    end else begin
      grt_wg_alloc_done <= _GEN_23;
    end
    if (reset) begin // @[top_resource_table.scala 136:38]
      grt_wg_dealloc_done <= 1'h0; // @[top_resource_table.scala 136:38]
    end else begin
      grt_wg_dealloc_done <= _GEN_24;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  done_array_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wf_count_array_0 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  wg_count_array_0 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  vgpr_start_array_0 = _RAND_3[12:0];
  _RAND_4 = {1{`RANDOM}};
  vgpr_size_array_0 = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  sgpr_start_array_0 = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  sgpr_size_array_0 = _RAND_6[12:0];
  _RAND_7 = {1{`RANDOM}};
  lds_start_array_0 = _RAND_7[12:0];
  _RAND_8 = {1{`RANDOM}};
  lds_size_array_0 = _RAND_8[12:0];
  _RAND_9 = {1{`RANDOM}};
  cu_id_array_0 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  serviced_array_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  is_alloc_array_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  done_cancelled_array_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  command_serviced_array_cancelled_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  grt_cam_up_valid_i = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  grt_wg_alloc_done = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  grt_wg_dealloc_done = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM(
  input         clock,
  input         reset,
  input         io_rd_addr,
  input         io_wr_addr,
  input  [57:0] io_wr_word,
  output [57:0] io_rd_word,
  input         io_wr_en,
  input         io_rd_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [57:0] mem [0:1]; // @[RAM.scala 14:18]
  wire  mem_rd_word_reg_MPORT_en; // @[RAM.scala 14:18]
  wire  mem_rd_word_reg_MPORT_addr; // @[RAM.scala 14:18]
  wire [57:0] mem_rd_word_reg_MPORT_data; // @[RAM.scala 14:18]
  wire [57:0] mem_MPORT_data; // @[RAM.scala 14:18]
  wire  mem_MPORT_addr; // @[RAM.scala 14:18]
  wire  mem_MPORT_mask; // @[RAM.scala 14:18]
  wire  mem_MPORT_en; // @[RAM.scala 14:18]
  reg [57:0] rd_word_reg; // @[RAM.scala 19:30]
  assign mem_rd_word_reg_MPORT_en = io_rd_en;
  assign mem_rd_word_reg_MPORT_addr = io_rd_addr;
  assign mem_rd_word_reg_MPORT_data = mem[mem_rd_word_reg_MPORT_addr]; // @[RAM.scala 14:18]
  assign mem_MPORT_data = io_wr_word;
  assign mem_MPORT_addr = io_wr_addr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wr_en;
  assign io_rd_word = rd_word_reg; // @[RAM.scala 23:16]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[RAM.scala 14:18]
    end
    if (reset) begin // @[RAM.scala 19:30]
      rd_word_reg <= 58'h0; // @[RAM.scala 19:30]
    end else if (io_rd_en) begin // @[RAM.scala 20:20]
      rd_word_reg <= mem_rd_word_reg_MPORT_data; // @[RAM.scala 21:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mem[initvar] = _RAND_0[57:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  rd_word_reg = _RAND_1[57:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_1(
  input         clock,
  input         reset,
  input         io_rd_addr,
  input         io_wr_addr,
  input  [72:0] io_wr_word,
  output [72:0] io_rd_word,
  input         io_wr_en,
  input         io_rd_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [72:0] mem [0:1]; // @[RAM.scala 14:18]
  wire  mem_rd_word_reg_MPORT_en; // @[RAM.scala 14:18]
  wire  mem_rd_word_reg_MPORT_addr; // @[RAM.scala 14:18]
  wire [72:0] mem_rd_word_reg_MPORT_data; // @[RAM.scala 14:18]
  wire [72:0] mem_MPORT_data; // @[RAM.scala 14:18]
  wire  mem_MPORT_addr; // @[RAM.scala 14:18]
  wire  mem_MPORT_mask; // @[RAM.scala 14:18]
  wire  mem_MPORT_en; // @[RAM.scala 14:18]
  reg [72:0] rd_word_reg; // @[RAM.scala 19:30]
  assign mem_rd_word_reg_MPORT_en = io_rd_en;
  assign mem_rd_word_reg_MPORT_addr = io_rd_addr;
  assign mem_rd_word_reg_MPORT_data = mem[mem_rd_word_reg_MPORT_addr]; // @[RAM.scala 14:18]
  assign mem_MPORT_data = io_wr_word;
  assign mem_MPORT_addr = io_wr_addr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wr_en;
  assign io_rd_word = rd_word_reg; // @[RAM.scala 23:16]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[RAM.scala 14:18]
    end
    if (reset) begin // @[RAM.scala 19:30]
      rd_word_reg <= 73'h0; // @[RAM.scala 19:30]
    end else if (io_rd_en) begin // @[RAM.scala 20:20]
      rd_word_reg <= mem_rd_word_reg_MPORT_data; // @[RAM.scala 21:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mem[initvar] = _RAND_0[72:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  rd_word_reg = _RAND_1[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module inflight_wg_buffer(
  input         clock,
  input         reset,
  input         io_host_wg_valid,
  input  [4:0]  io_host_wg_id,
  input  [2:0]  io_host_num_wf,
  input  [9:0]  io_host_wf_size,
  input  [31:0] io_host_start_pc,
  input  [12:0] io_host_vgpr_size_total,
  input  [12:0] io_host_sgpr_size_total,
  input  [12:0] io_host_lds_size_total,
  input  [10:0] io_host_gds_size_total,
  input  [12:0] io_host_vgpr_size_per_wf,
  input  [12:0] io_host_sgpr_size_per_wf,
  input         io_dis_controller_wg_alloc_valid,
  input         io_dis_controller_start_alloc,
  input         io_dis_controller_wg_dealloc_valid,
  input         io_dis_controller_wg_rejected_valid,
  input  [4:0]  io_allocator_wg_id_out,
  input  [4:0]  io_gpu_interface_dealloc_wg_id,
  output        io_inflight_wg_buffer_host_rcvd_ack,
  output        io_inflight_wg_buffer_host_wf_done,
  output [4:0]  io_inflight_wg_buffer_host_wf_done_wg_id,
  output        io_inflight_wg_buffer_alloc_valid,
  output        io_inflight_wg_buffer_alloc_available,
  output [4:0]  io_inflight_wg_buffer_alloc_wg_id,
  output [2:0]  io_inflight_wg_buffer_alloc_num_wf,
  output [12:0] io_inflight_wg_buffer_alloc_vgpr_size,
  output [12:0] io_inflight_wg_buffer_alloc_sgpr_size,
  output [12:0] io_inflight_wg_buffer_alloc_lds_size,
  output        io_inflight_wg_buffer_gpu_valid,
  output [12:0] io_inflight_wg_buffer_gpu_vgpr_size_per_wf,
  output [12:0] io_inflight_wg_buffer_gpu_sgpr_size_per_wf,
  output [9:0]  io_inflight_wg_buffer_gpu_wf_size,
  output [31:0] io_inflight_wg_buffer_start_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [95:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  wire  ram_wg_waiting_allocation_clock; // @[inflight_wg_buffer.scala 94:43]
  wire  ram_wg_waiting_allocation_reset; // @[inflight_wg_buffer.scala 94:43]
  wire  ram_wg_waiting_allocation_io_rd_addr; // @[inflight_wg_buffer.scala 94:43]
  wire  ram_wg_waiting_allocation_io_wr_addr; // @[inflight_wg_buffer.scala 94:43]
  wire [57:0] ram_wg_waiting_allocation_io_wr_word; // @[inflight_wg_buffer.scala 94:43]
  wire [57:0] ram_wg_waiting_allocation_io_rd_word; // @[inflight_wg_buffer.scala 94:43]
  wire  ram_wg_waiting_allocation_io_wr_en; // @[inflight_wg_buffer.scala 94:43]
  wire  ram_wg_waiting_allocation_io_rd_en; // @[inflight_wg_buffer.scala 94:43]
  wire  ram_wg_ready_start_clock; // @[inflight_wg_buffer.scala 98:36]
  wire  ram_wg_ready_start_reset; // @[inflight_wg_buffer.scala 98:36]
  wire  ram_wg_ready_start_io_rd_addr; // @[inflight_wg_buffer.scala 98:36]
  wire  ram_wg_ready_start_io_wr_addr; // @[inflight_wg_buffer.scala 98:36]
  wire [72:0] ram_wg_ready_start_io_wr_word; // @[inflight_wg_buffer.scala 98:36]
  wire [72:0] ram_wg_ready_start_io_rd_word; // @[inflight_wg_buffer.scala 98:36]
  wire  ram_wg_ready_start_io_wr_en; // @[inflight_wg_buffer.scala 98:36]
  wire  ram_wg_ready_start_io_rd_en; // @[inflight_wg_buffer.scala 98:36]
  reg  host_wg_valid_i; // @[inflight_wg_buffer.scala 131:34]
  reg [4:0] host_wg_id_i; // @[inflight_wg_buffer.scala 133:31]
  reg [2:0] host_num_wf_i; // @[inflight_wg_buffer.scala 135:32]
  reg [9:0] host_wf_size_i; // @[inflight_wg_buffer.scala 137:33]
  reg [31:0] host_start_pc_i; // @[inflight_wg_buffer.scala 139:34]
  reg [12:0] host_vgpr_size_total_i; // @[inflight_wg_buffer.scala 141:41]
  reg [12:0] host_sgpr_size_total_i; // @[inflight_wg_buffer.scala 143:41]
  reg [12:0] host_vgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 145:42]
  reg [12:0] host_sgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 147:42]
  reg [12:0] host_lds_size_total_i; // @[inflight_wg_buffer.scala 149:40]
  reg [10:0] host_gds_size_total_i; // @[inflight_wg_buffer.scala 151:40]
  reg  dis_controller_start_alloc_i; // @[inflight_wg_buffer.scala 153:47]
  reg  dis_controller_wg_alloc_valid_i; // @[inflight_wg_buffer.scala 155:50]
  reg  dis_controller_wg_dealloc_valid_i; // @[inflight_wg_buffer.scala 156:52]
  reg  dis_controller_wg_rejected_valid_i; // @[inflight_wg_buffer.scala 157:53]
  reg [4:0] gpu_interface_dealloc_wg_id_i; // @[inflight_wg_buffer.scala 160:48]
  reg [7:0] inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 162:40]
  reg [3:0] inflight_tbl_rd_host_st; // @[inflight_wg_buffer.scala 163:42]
  reg [4:0] allocator_wg_id_out_i; // @[inflight_wg_buffer.scala 164:40]
  wire  _GEN_0 = io_dis_controller_wg_alloc_valid | dis_controller_wg_alloc_valid_i; // @[inflight_wg_buffer.scala 165:43 166:39 155:50]
  wire  _GEN_2 = io_dis_controller_wg_rejected_valid | dis_controller_wg_rejected_valid_i; // @[inflight_wg_buffer.scala 169:46 170:42 157:53]
  reg  inflight_wg_buffer_host_wf_done_i; // @[inflight_wg_buffer.scala 173:52]
  reg [4:0] inflight_wg_buffer_host_wf_done_wg_id_i; // @[inflight_wg_buffer.scala 175:58]
  reg  waiting_tbl_valid_0; // @[inflight_wg_buffer.scala 185:36]
  reg  waiting_tbl_valid_1; // @[inflight_wg_buffer.scala 185:36]
  reg  new_index_wr_en; // @[inflight_wg_buffer.scala 186:34]
  reg [57:0] new_entry_wg_reg; // @[inflight_wg_buffer.scala 189:35]
  reg [72:0] ready_tbl_wr_reg; // @[inflight_wg_buffer.scala 191:35]
  reg  inflight_wg_buffer_host_rcvd_ack_i; // @[inflight_wg_buffer.scala 193:53]
  reg  new_index; // @[inflight_wg_buffer.scala 195:28]
  wire  _T_1 = ~waiting_tbl_valid_0; // @[inflight_wg_buffer.scala 212:42]
  wire  _T_2 = ~waiting_tbl_valid_1; // @[inflight_wg_buffer.scala 212:42]
  wire [57:0] _new_entry_wg_reg_T = {host_num_wf_i,host_lds_size_total_i,host_gds_size_total_i,host_wg_id_i,
    host_vgpr_size_total_i,host_sgpr_size_total_i}; // @[Cat.scala 31:58]
  wire [72:0] _ready_tbl_wr_reg_T = {host_start_pc_i,host_wf_size_i,host_wg_id_i,host_vgpr_size_per_wf_i,
    host_sgpr_size_per_wf_i}; // @[Cat.scala 31:58]
  wire  _GEN_8 = ~new_index | waiting_tbl_valid_0; // @[inflight_wg_buffer.scala 185:36 233:{38,38}]
  wire  _GEN_9 = new_index | waiting_tbl_valid_1; // @[inflight_wg_buffer.scala 185:36 233:{38,38}]
  wire [3:0] _GEN_10 = 4'h8 == inflight_tbl_rd_host_st ? 4'h1 : inflight_tbl_rd_host_st; // @[inflight_wg_buffer.scala 205:36 240:33 163:42]
  wire  _GEN_11 = 4'h4 == inflight_tbl_rd_host_st ? _GEN_8 : waiting_tbl_valid_0; // @[inflight_wg_buffer.scala 185:36 205:36]
  wire  _GEN_12 = 4'h4 == inflight_tbl_rd_host_st ? _GEN_9 : waiting_tbl_valid_1; // @[inflight_wg_buffer.scala 185:36 205:36]
  wire  _GEN_18 = 4'h2 == inflight_tbl_rd_host_st ? waiting_tbl_valid_0 : _GEN_11; // @[inflight_wg_buffer.scala 185:36 205:36]
  wire  _GEN_19 = 4'h2 == inflight_tbl_rd_host_st ? waiting_tbl_valid_1 : _GEN_12; // @[inflight_wg_buffer.scala 185:36 205:36]
  wire  _GEN_24 = 4'h1 == inflight_tbl_rd_host_st ? waiting_tbl_valid_0 : _GEN_18; // @[inflight_wg_buffer.scala 185:36 205:36]
  wire  _GEN_25 = 4'h1 == inflight_tbl_rd_host_st ? waiting_tbl_valid_1 : _GEN_19; // @[inflight_wg_buffer.scala 185:36 205:36]
  reg  waiting_tbl_pending_0; // @[inflight_wg_buffer.scala 245:38]
  reg  waiting_tbl_pending_1; // @[inflight_wg_buffer.scala 245:38]
  reg  chosen_entry; // @[inflight_wg_buffer.scala 246:31]
  reg  chosen_entry_by_allocator; // @[inflight_wg_buffer.scala 247:44]
  reg  chosen_entry_is_valid; // @[inflight_wg_buffer.scala 248:40]
  reg  wait_tbl_busy; // @[inflight_wg_buffer.scala 249:32]
  wire  valid_not_pending_0 = waiting_tbl_valid_0 & ~waiting_tbl_pending_0; // @[inflight_wg_buffer.scala 254:52]
  wire  valid_not_pending_1 = waiting_tbl_valid_1 & ~waiting_tbl_pending_1; // @[inflight_wg_buffer.scala 254:52]
  reg [4:0] tbl_walk_wg_id_searched; // @[inflight_wg_buffer.scala 257:42]
  reg  tbl_walk_rd_en; // @[inflight_wg_buffer.scala 262:33]
  reg  tbl_walk_idx; // @[inflight_wg_buffer.scala 265:31]
  reg  tbl_walk_rd_valid; // @[inflight_wg_buffer.scala 268:36]
  reg  inflight_wg_buffer_gpu_valid_i; // @[inflight_wg_buffer.scala 274:49]
  reg [12:0] inflight_wg_buffer_gpu_vgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 276:60]
  reg [12:0] inflight_wg_buffer_gpu_sgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 278:60]
  reg [9:0] inflight_wg_buffer_gpu_wf_size_i; // @[inflight_wg_buffer.scala 280:51]
  reg [31:0] inflight_wg_buffer_start_pc_i; // @[inflight_wg_buffer.scala 282:48]
  reg [4:0] inflight_wg_buffer_alloc_wg_id_i; // @[inflight_wg_buffer.scala 286:51]
  reg [2:0] inflight_wg_buffer_alloc_num_wf_i; // @[inflight_wg_buffer.scala 288:52]
  reg [12:0] inflight_wg_buffer_alloc_vgpr_size_i; // @[inflight_wg_buffer.scala 290:55]
  reg [12:0] inflight_wg_buffer_alloc_sgpr_size_i; // @[inflight_wg_buffer.scala 292:55]
  reg [12:0] inflight_wg_buffer_alloc_lds_size_i; // @[inflight_wg_buffer.scala 294:54]
  reg  wg_waiting_alloc_valid; // @[inflight_wg_buffer.scala 298:41]
  reg  last_chosen_entry_rr; // @[inflight_wg_buffer.scala 300:39]
  wire  _GEN_26 = dis_controller_start_alloc_i ? chosen_entry_by_allocator : last_chosen_entry_rr; // @[inflight_wg_buffer.scala 301:39 302:28 300:39]
  wire  _GEN_27 = ~chosen_entry_by_allocator | waiting_tbl_pending_0; // @[inflight_wg_buffer.scala 245:38 313:{58,58}]
  wire  _GEN_28 = chosen_entry_by_allocator | waiting_tbl_pending_1; // @[inflight_wg_buffer.scala 245:38 313:{58,58}]
  wire  _T_14 = ~wg_waiting_alloc_valid & (valid_not_pending_0 | valid_not_pending_1); // @[inflight_wg_buffer.scala 317:43]
  wire  _GEN_35 = dis_controller_start_alloc_i | _T_14; // @[inflight_wg_buffer.scala 250:19 312:43]
  wire  _GEN_36 = dis_controller_wg_rejected_valid_i ? 1'h0 : _GEN_2; // @[inflight_wg_buffer.scala 339:54 340:46]
  wire [4:0] _GEN_37 = dis_controller_wg_rejected_valid_i ? allocator_wg_id_out_i : tbl_walk_wg_id_searched; // @[inflight_wg_buffer.scala 339:54 341:35 257:42]
  wire  _GEN_39 = dis_controller_wg_rejected_valid_i ? 1'h0 : tbl_walk_idx; // @[inflight_wg_buffer.scala 339:54 344:24 265:31]
  wire [7:0] _GEN_40 = dis_controller_wg_rejected_valid_i ? 8'h10 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 339:54 345:33 162:40]
  wire  _GEN_43 = dis_controller_wg_alloc_valid_i | dis_controller_wg_rejected_valid_i; // @[inflight_wg_buffer.scala 330:46 333:26]
  wire [57:0] table_walk_rd_reg = ram_wg_waiting_allocation_io_rd_word; // @[inflight_wg_buffer.scala 258:33 259:23]
  wire  _GEN_48 = tbl_walk_idx ? waiting_tbl_pending_1 : waiting_tbl_pending_0; // @[inflight_wg_buffer.scala 354:{82,82}]
  wire  _T_19 = table_walk_rd_reg[30:26] == tbl_walk_wg_id_searched & _GEN_48; // @[inflight_wg_buffer.scala 354:82]
  wire [7:0] _GEN_49 = table_walk_rd_reg[30:26] == tbl_walk_wg_id_searched & _GEN_48 ? 8'h8 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 354:119 356:35 162:40]
  wire  _GEN_50 = table_walk_rd_reg[30:26] == tbl_walk_wg_id_searched & _GEN_48 ? tbl_walk_idx : tbl_walk_idx + 1'h1; // @[inflight_wg_buffer.scala 354:119 265:31 359:26]
  wire  _GEN_51 = table_walk_rd_reg[30:26] == tbl_walk_wg_id_searched & _GEN_48 ? 1'h0 : 1'h1; // @[inflight_wg_buffer.scala 354:119 271:20 360:28]
  wire [7:0] _GEN_52 = tbl_walk_rd_valid ? _GEN_49 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 353:32 162:40]
  wire  _GEN_53 = tbl_walk_rd_valid ? _GEN_50 : tbl_walk_idx; // @[inflight_wg_buffer.scala 265:31 353:32]
  wire  _GEN_54 = tbl_walk_rd_valid & _GEN_51; // @[inflight_wg_buffer.scala 271:20 353:32]
  wire  _GEN_55 = ~tbl_walk_idx ? 1'h0 : _GEN_24; // @[inflight_wg_buffer.scala 366:{41,41}]
  wire  _GEN_56 = tbl_walk_idx ? 1'h0 : _GEN_25; // @[inflight_wg_buffer.scala 366:{41,41}]
  wire  _GEN_57 = ~tbl_walk_idx ? 1'h0 : waiting_tbl_pending_0; // @[inflight_wg_buffer.scala 245:38 367:{43,43}]
  wire  _GEN_58 = tbl_walk_idx ? 1'h0 : waiting_tbl_pending_1; // @[inflight_wg_buffer.scala 245:38 367:{43,43}]
  wire [72:0] ready_tbl_rd_reg = ram_wg_ready_start_io_rd_word; // @[inflight_wg_buffer.scala 260:32 261:22]
  wire [7:0] _GEN_59 = _T_19 ? 8'h20 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 381:119 382:35 162:40]
  wire [7:0] _GEN_62 = tbl_walk_rd_valid ? _GEN_59 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 380:32 162:40]
  wire  _GEN_68 = chosen_entry_is_valid ? chosen_entry : tbl_walk_idx; // @[inflight_wg_buffer.scala 399:36 401:24 265:31]
  wire  _GEN_69 = chosen_entry_is_valid ? chosen_entry : chosen_entry_by_allocator; // @[inflight_wg_buffer.scala 399:36 402:37 247:44]
  wire [7:0] _GEN_70 = chosen_entry_is_valid ? 8'h80 : 8'h1; // @[inflight_wg_buffer.scala 399:36 403:33 406:33]
  wire  _GEN_71 = tbl_walk_rd_valid | wg_waiting_alloc_valid; // @[inflight_wg_buffer.scala 413:32 414:34 298:41]
  wire [4:0] _GEN_72 = tbl_walk_rd_valid ? table_walk_rd_reg[30:26] : inflight_wg_buffer_alloc_wg_id_i; // @[inflight_wg_buffer.scala 413:32 415:44 286:51]
  wire [2:0] _GEN_73 = tbl_walk_rd_valid ? table_walk_rd_reg[57:55] : inflight_wg_buffer_alloc_num_wf_i; // @[inflight_wg_buffer.scala 413:32 416:45 288:52]
  wire [12:0] _GEN_74 = tbl_walk_rd_valid ? table_walk_rd_reg[25:13] : inflight_wg_buffer_alloc_vgpr_size_i; // @[inflight_wg_buffer.scala 413:32 417:48 290:55]
  wire [12:0] _GEN_75 = tbl_walk_rd_valid ? table_walk_rd_reg[12:0] : inflight_wg_buffer_alloc_sgpr_size_i; // @[inflight_wg_buffer.scala 413:32 418:48 292:55]
  wire [12:0] _GEN_76 = tbl_walk_rd_valid ? table_walk_rd_reg[54:42] : inflight_wg_buffer_alloc_lds_size_i; // @[inflight_wg_buffer.scala 413:32 419:47 294:54]
  wire [7:0] _GEN_78 = tbl_walk_rd_valid ? 8'h1 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 413:32 421:33 162:40]
  wire  _GEN_79 = 8'h80 == inflight_tbl_alloc_st ? _GEN_71 : wg_waiting_alloc_valid; // @[inflight_wg_buffer.scala 306:34 298:41]
  wire [4:0] _GEN_80 = 8'h80 == inflight_tbl_alloc_st ? _GEN_72 : inflight_wg_buffer_alloc_wg_id_i; // @[inflight_wg_buffer.scala 306:34 286:51]
  wire [2:0] _GEN_81 = 8'h80 == inflight_tbl_alloc_st ? _GEN_73 : inflight_wg_buffer_alloc_num_wf_i; // @[inflight_wg_buffer.scala 306:34 288:52]
  wire [12:0] _GEN_82 = 8'h80 == inflight_tbl_alloc_st ? _GEN_74 : inflight_wg_buffer_alloc_vgpr_size_i; // @[inflight_wg_buffer.scala 306:34 290:55]
  wire [12:0] _GEN_83 = 8'h80 == inflight_tbl_alloc_st ? _GEN_75 : inflight_wg_buffer_alloc_sgpr_size_i; // @[inflight_wg_buffer.scala 306:34 292:55]
  wire [12:0] _GEN_84 = 8'h80 == inflight_tbl_alloc_st ? _GEN_76 : inflight_wg_buffer_alloc_lds_size_i; // @[inflight_wg_buffer.scala 306:34 294:54]
  wire [7:0] _GEN_86 = 8'h80 == inflight_tbl_alloc_st ? _GEN_78 : inflight_tbl_alloc_st; // @[inflight_wg_buffer.scala 306:34 162:40]
  wire  _GEN_88 = 8'h40 == inflight_tbl_alloc_st ? _GEN_68 : tbl_walk_idx; // @[inflight_wg_buffer.scala 265:31 306:34]
  wire  _GEN_89 = 8'h40 == inflight_tbl_alloc_st ? _GEN_69 : chosen_entry_by_allocator; // @[inflight_wg_buffer.scala 306:34 247:44]
  wire [7:0] _GEN_90 = 8'h40 == inflight_tbl_alloc_st ? _GEN_70 : _GEN_86; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_91 = 8'h40 == inflight_tbl_alloc_st ? wg_waiting_alloc_valid : _GEN_79; // @[inflight_wg_buffer.scala 306:34 298:41]
  wire [4:0] _GEN_92 = 8'h40 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_wg_id_i : _GEN_80; // @[inflight_wg_buffer.scala 306:34 286:51]
  wire [2:0] _GEN_93 = 8'h40 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_num_wf_i : _GEN_81; // @[inflight_wg_buffer.scala 306:34 288:52]
  wire [12:0] _GEN_94 = 8'h40 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_vgpr_size_i : _GEN_82; // @[inflight_wg_buffer.scala 306:34 290:55]
  wire [12:0] _GEN_95 = 8'h40 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_sgpr_size_i : _GEN_83; // @[inflight_wg_buffer.scala 306:34 292:55]
  wire [12:0] _GEN_96 = 8'h40 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_lds_size_i : _GEN_84; // @[inflight_wg_buffer.scala 306:34 294:54]
  wire  _GEN_98 = 8'h20 == inflight_tbl_alloc_st ? _GEN_57 : waiting_tbl_pending_0; // @[inflight_wg_buffer.scala 306:34 245:38]
  wire  _GEN_99 = 8'h20 == inflight_tbl_alloc_st ? _GEN_58 : waiting_tbl_pending_1; // @[inflight_wg_buffer.scala 306:34 245:38]
  wire [7:0] _GEN_100 = 8'h20 == inflight_tbl_alloc_st ? 8'h40 : _GEN_90; // @[inflight_wg_buffer.scala 306:34 392:31]
  wire  _GEN_101 = 8'h20 == inflight_tbl_alloc_st ? 1'h0 : 8'h40 == inflight_tbl_alloc_st & chosen_entry_is_valid; // @[inflight_wg_buffer.scala 271:20 306:34]
  wire  _GEN_102 = 8'h20 == inflight_tbl_alloc_st ? tbl_walk_idx : _GEN_88; // @[inflight_wg_buffer.scala 265:31 306:34]
  wire  _GEN_103 = 8'h20 == inflight_tbl_alloc_st ? chosen_entry_by_allocator : _GEN_89; // @[inflight_wg_buffer.scala 306:34 247:44]
  wire  _GEN_104 = 8'h20 == inflight_tbl_alloc_st ? wg_waiting_alloc_valid : _GEN_91; // @[inflight_wg_buffer.scala 306:34 298:41]
  wire [4:0] _GEN_105 = 8'h20 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_wg_id_i : _GEN_92; // @[inflight_wg_buffer.scala 306:34 286:51]
  wire [2:0] _GEN_106 = 8'h20 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_num_wf_i : _GEN_93; // @[inflight_wg_buffer.scala 306:34 288:52]
  wire [12:0] _GEN_107 = 8'h20 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_vgpr_size_i : _GEN_94; // @[inflight_wg_buffer.scala 306:34 290:55]
  wire [12:0] _GEN_108 = 8'h20 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_sgpr_size_i : _GEN_95; // @[inflight_wg_buffer.scala 306:34 292:55]
  wire [12:0] _GEN_109 = 8'h20 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_lds_size_i : _GEN_96; // @[inflight_wg_buffer.scala 306:34 294:54]
  wire [7:0] _GEN_111 = 8'h10 == inflight_tbl_alloc_st ? _GEN_62 : _GEN_100; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_112 = 8'h10 == inflight_tbl_alloc_st ? _GEN_53 : _GEN_102; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_113 = 8'h10 == inflight_tbl_alloc_st ? _GEN_54 : _GEN_101; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_114 = 8'h10 == inflight_tbl_alloc_st ? waiting_tbl_pending_0 : _GEN_98; // @[inflight_wg_buffer.scala 306:34 245:38]
  wire  _GEN_115 = 8'h10 == inflight_tbl_alloc_st ? waiting_tbl_pending_1 : _GEN_99; // @[inflight_wg_buffer.scala 306:34 245:38]
  wire  _GEN_116 = 8'h10 == inflight_tbl_alloc_st ? chosen_entry_by_allocator : _GEN_103; // @[inflight_wg_buffer.scala 306:34 247:44]
  wire  _GEN_117 = 8'h10 == inflight_tbl_alloc_st ? wg_waiting_alloc_valid : _GEN_104; // @[inflight_wg_buffer.scala 306:34 298:41]
  wire [4:0] _GEN_118 = 8'h10 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_wg_id_i : _GEN_105; // @[inflight_wg_buffer.scala 306:34 286:51]
  wire [2:0] _GEN_119 = 8'h10 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_num_wf_i : _GEN_106; // @[inflight_wg_buffer.scala 306:34 288:52]
  wire [12:0] _GEN_120 = 8'h10 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_vgpr_size_i : _GEN_107; // @[inflight_wg_buffer.scala 306:34 290:55]
  wire [12:0] _GEN_121 = 8'h10 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_sgpr_size_i : _GEN_108; // @[inflight_wg_buffer.scala 306:34 292:55]
  wire [12:0] _GEN_122 = 8'h10 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_lds_size_i : _GEN_109; // @[inflight_wg_buffer.scala 306:34 294:54]
  wire  _GEN_124 = 8'h8 == inflight_tbl_alloc_st ? _GEN_55 : _GEN_24; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_125 = 8'h8 == inflight_tbl_alloc_st ? _GEN_56 : _GEN_25; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_126 = 8'h8 == inflight_tbl_alloc_st ? _GEN_57 : _GEN_114; // @[inflight_wg_buffer.scala 306:34]
  wire  _GEN_127 = 8'h8 == inflight_tbl_alloc_st ? _GEN_58 : _GEN_115; // @[inflight_wg_buffer.scala 306:34]
  wire [12:0] _GEN_129 = 8'h8 == inflight_tbl_alloc_st ? ready_tbl_rd_reg[25:13] :
    inflight_wg_buffer_gpu_vgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 306:34 369:51 276:60]
  wire [12:0] _GEN_130 = 8'h8 == inflight_tbl_alloc_st ? ready_tbl_rd_reg[12:0] :
    inflight_wg_buffer_gpu_sgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 306:34 370:51 278:60]
  wire [9:0] _GEN_131 = 8'h8 == inflight_tbl_alloc_st ? ready_tbl_rd_reg[40:31] : inflight_wg_buffer_gpu_wf_size_i; // @[inflight_wg_buffer.scala 306:34 371:42 280:51]
  wire [31:0] _GEN_132 = 8'h8 == inflight_tbl_alloc_st ? ready_tbl_rd_reg[72:41] : inflight_wg_buffer_start_pc_i; // @[inflight_wg_buffer.scala 306:34 372:39 282:48]
  wire [7:0] _GEN_133 = 8'h8 == inflight_tbl_alloc_st ? 8'h40 : _GEN_111; // @[inflight_wg_buffer.scala 306:34 373:31]
  wire  _GEN_134 = 8'h8 == inflight_tbl_alloc_st ? tbl_walk_idx : _GEN_112; // @[inflight_wg_buffer.scala 265:31 306:34]
  wire  _GEN_135 = 8'h8 == inflight_tbl_alloc_st ? 1'h0 : _GEN_113; // @[inflight_wg_buffer.scala 271:20 306:34]
  wire  _GEN_136 = 8'h8 == inflight_tbl_alloc_st ? chosen_entry_by_allocator : _GEN_116; // @[inflight_wg_buffer.scala 306:34 247:44]
  wire  _GEN_137 = 8'h8 == inflight_tbl_alloc_st ? wg_waiting_alloc_valid : _GEN_117; // @[inflight_wg_buffer.scala 306:34 298:41]
  wire [4:0] _GEN_138 = 8'h8 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_wg_id_i : _GEN_118; // @[inflight_wg_buffer.scala 306:34 286:51]
  wire [2:0] _GEN_139 = 8'h8 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_num_wf_i : _GEN_119; // @[inflight_wg_buffer.scala 306:34 288:52]
  wire [12:0] _GEN_140 = 8'h8 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_vgpr_size_i : _GEN_120; // @[inflight_wg_buffer.scala 306:34 290:55]
  wire [12:0] _GEN_141 = 8'h8 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_sgpr_size_i : _GEN_121; // @[inflight_wg_buffer.scala 306:34 292:55]
  wire [12:0] _GEN_142 = 8'h8 == inflight_tbl_alloc_st ? inflight_wg_buffer_alloc_lds_size_i : _GEN_122; // @[inflight_wg_buffer.scala 306:34 294:54]
  wire  _left_degree_T_1 = 1'h1 + last_chosen_entry_rr; // @[inflight_wg_buffer.scala 449:56]
  wire [1:0] _GEN_231 = {{1'd0}, _left_degree_T_1}; // @[inflight_wg_buffer.scala 449:49]
  wire [1:0] left_degree = 2'h2 - _GEN_231; // @[inflight_wg_buffer.scala 449:49]
  wire [1:0] _waiting_tbl_valid_rotated_0_T_1 = 2'h0 - left_degree; // @[inflight_wg_buffer.scala 453:63]
  wire  _GEN_216 = _waiting_tbl_valid_rotated_0_T_1[0] ? valid_not_pending_1 : valid_not_pending_0; // @[inflight_wg_buffer.scala 453:{38,38}]
  wire  _GEN_218 = _GEN_231[0] ? valid_not_pending_1 : valid_not_pending_0; // @[inflight_wg_buffer.scala 456:{38,38}]
  wire  waiting_tbl_valid_rotated_0 = 2'h0 >= left_degree ? _GEN_216 : _GEN_218; // @[inflight_wg_buffer.scala 452:31 453:38 456:38]
  wire [1:0] _waiting_tbl_valid_rotated_1_T_1 = 2'h1 - left_degree; // @[inflight_wg_buffer.scala 453:63]
  wire  _GEN_221 = _waiting_tbl_valid_rotated_1_T_1[0] ? valid_not_pending_1 : valid_not_pending_0; // @[inflight_wg_buffer.scala 453:{38,38}]
  wire  _GEN_223 = 1'h1 + _left_degree_T_1 ? valid_not_pending_1 : valid_not_pending_0; // @[inflight_wg_buffer.scala 456:{38,38}]
  wire  waiting_tbl_valid_rotated_1 = 2'h1 >= left_degree ? _GEN_221 : _GEN_223; // @[inflight_wg_buffer.scala 452:31 453:38 456:38]
  wire  _GEN_226 = waiting_tbl_valid_rotated_1 & _left_degree_T_1 + 1'h1; // @[inflight_wg_buffer.scala 448:23 460:41 462:27]
  wire [1:0] _idx_found_entry_c_T_4 = {{1'd0}, last_chosen_entry_rr}; // @[inflight_wg_buffer.scala 462:34]
  wire  found_entry_valid_c = waiting_tbl_valid_rotated_0 | waiting_tbl_valid_rotated_1; // @[inflight_wg_buffer.scala 460:41 461:29]
  RAM ram_wg_waiting_allocation ( // @[inflight_wg_buffer.scala 94:43]
    .clock(ram_wg_waiting_allocation_clock),
    .reset(ram_wg_waiting_allocation_reset),
    .io_rd_addr(ram_wg_waiting_allocation_io_rd_addr),
    .io_wr_addr(ram_wg_waiting_allocation_io_wr_addr),
    .io_wr_word(ram_wg_waiting_allocation_io_wr_word),
    .io_rd_word(ram_wg_waiting_allocation_io_rd_word),
    .io_wr_en(ram_wg_waiting_allocation_io_wr_en),
    .io_rd_en(ram_wg_waiting_allocation_io_rd_en)
  );
  RAM_1 ram_wg_ready_start ( // @[inflight_wg_buffer.scala 98:36]
    .clock(ram_wg_ready_start_clock),
    .reset(ram_wg_ready_start_reset),
    .io_rd_addr(ram_wg_ready_start_io_rd_addr),
    .io_wr_addr(ram_wg_ready_start_io_wr_addr),
    .io_wr_word(ram_wg_ready_start_io_wr_word),
    .io_rd_word(ram_wg_ready_start_io_rd_word),
    .io_wr_en(ram_wg_ready_start_io_wr_en),
    .io_rd_en(ram_wg_ready_start_io_rd_en)
  );
  assign io_inflight_wg_buffer_host_rcvd_ack = inflight_wg_buffer_host_rcvd_ack_i; // @[inflight_wg_buffer.scala 194:41]
  assign io_inflight_wg_buffer_host_wf_done = inflight_wg_buffer_host_wf_done_i; // @[inflight_wg_buffer.scala 174:40]
  assign io_inflight_wg_buffer_host_wf_done_wg_id = inflight_wg_buffer_host_wf_done_wg_id_i; // @[inflight_wg_buffer.scala 176:46]
  assign io_inflight_wg_buffer_alloc_valid = wg_waiting_alloc_valid; // @[inflight_wg_buffer.scala 299:39]
  assign io_inflight_wg_buffer_alloc_available = ~wait_tbl_busy; // @[inflight_wg_buffer.scala 251:46]
  assign io_inflight_wg_buffer_alloc_wg_id = inflight_wg_buffer_alloc_wg_id_i; // @[inflight_wg_buffer.scala 287:39]
  assign io_inflight_wg_buffer_alloc_num_wf = inflight_wg_buffer_alloc_num_wf_i; // @[inflight_wg_buffer.scala 289:40]
  assign io_inflight_wg_buffer_alloc_vgpr_size = inflight_wg_buffer_alloc_vgpr_size_i; // @[inflight_wg_buffer.scala 291:43]
  assign io_inflight_wg_buffer_alloc_sgpr_size = inflight_wg_buffer_alloc_sgpr_size_i; // @[inflight_wg_buffer.scala 293:43]
  assign io_inflight_wg_buffer_alloc_lds_size = inflight_wg_buffer_alloc_lds_size_i; // @[inflight_wg_buffer.scala 295:42]
  assign io_inflight_wg_buffer_gpu_valid = inflight_wg_buffer_gpu_valid_i; // @[inflight_wg_buffer.scala 275:37]
  assign io_inflight_wg_buffer_gpu_vgpr_size_per_wf = inflight_wg_buffer_gpu_vgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 277:48]
  assign io_inflight_wg_buffer_gpu_sgpr_size_per_wf = inflight_wg_buffer_gpu_sgpr_size_per_wf_i; // @[inflight_wg_buffer.scala 279:48]
  assign io_inflight_wg_buffer_gpu_wf_size = inflight_wg_buffer_gpu_wf_size_i; // @[inflight_wg_buffer.scala 281:39]
  assign io_inflight_wg_buffer_start_pc = inflight_wg_buffer_start_pc_i; // @[inflight_wg_buffer.scala 283:36]
  assign ram_wg_waiting_allocation_clock = clock;
  assign ram_wg_waiting_allocation_reset = reset;
  assign ram_wg_waiting_allocation_io_rd_addr = tbl_walk_idx; // @[inflight_wg_buffer.scala 266:42]
  assign ram_wg_waiting_allocation_io_wr_addr = new_index; // @[inflight_wg_buffer.scala 196:42]
  assign ram_wg_waiting_allocation_io_wr_word = new_entry_wg_reg; // @[inflight_wg_buffer.scala 190:42]
  assign ram_wg_waiting_allocation_io_wr_en = new_index_wr_en; // @[inflight_wg_buffer.scala 187:40]
  assign ram_wg_waiting_allocation_io_rd_en = tbl_walk_rd_en; // @[inflight_wg_buffer.scala 263:40]
  assign ram_wg_ready_start_clock = clock;
  assign ram_wg_ready_start_reset = reset;
  assign ram_wg_ready_start_io_rd_addr = tbl_walk_idx; // @[inflight_wg_buffer.scala 267:35]
  assign ram_wg_ready_start_io_wr_addr = new_index; // @[inflight_wg_buffer.scala 197:35]
  assign ram_wg_ready_start_io_wr_word = ready_tbl_wr_reg; // @[inflight_wg_buffer.scala 192:35]
  assign ram_wg_ready_start_io_wr_en = new_index_wr_en; // @[inflight_wg_buffer.scala 188:33]
  assign ram_wg_ready_start_io_rd_en = tbl_walk_rd_en; // @[inflight_wg_buffer.scala 264:33]
  always @(posedge clock) begin
    if (reset) begin // @[inflight_wg_buffer.scala 131:34]
      host_wg_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 131:34]
    end else begin
      host_wg_valid_i <= io_host_wg_valid; // @[inflight_wg_buffer.scala 132:21]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 133:31]
      host_wg_id_i <= 5'h0; // @[inflight_wg_buffer.scala 133:31]
    end else begin
      host_wg_id_i <= io_host_wg_id; // @[inflight_wg_buffer.scala 134:18]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 135:32]
      host_num_wf_i <= 3'h0; // @[inflight_wg_buffer.scala 135:32]
    end else begin
      host_num_wf_i <= io_host_num_wf; // @[inflight_wg_buffer.scala 136:19]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 137:33]
      host_wf_size_i <= 10'h0; // @[inflight_wg_buffer.scala 137:33]
    end else begin
      host_wf_size_i <= io_host_wf_size; // @[inflight_wg_buffer.scala 138:20]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 139:34]
      host_start_pc_i <= 32'h0; // @[inflight_wg_buffer.scala 139:34]
    end else begin
      host_start_pc_i <= io_host_start_pc; // @[inflight_wg_buffer.scala 140:21]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 141:41]
      host_vgpr_size_total_i <= 13'h0; // @[inflight_wg_buffer.scala 141:41]
    end else begin
      host_vgpr_size_total_i <= io_host_vgpr_size_total; // @[inflight_wg_buffer.scala 142:28]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 143:41]
      host_sgpr_size_total_i <= 13'h0; // @[inflight_wg_buffer.scala 143:41]
    end else begin
      host_sgpr_size_total_i <= io_host_sgpr_size_total; // @[inflight_wg_buffer.scala 144:28]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 145:42]
      host_vgpr_size_per_wf_i <= 13'h0; // @[inflight_wg_buffer.scala 145:42]
    end else begin
      host_vgpr_size_per_wf_i <= io_host_vgpr_size_per_wf; // @[inflight_wg_buffer.scala 146:29]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 147:42]
      host_sgpr_size_per_wf_i <= 13'h0; // @[inflight_wg_buffer.scala 147:42]
    end else begin
      host_sgpr_size_per_wf_i <= io_host_sgpr_size_per_wf; // @[inflight_wg_buffer.scala 148:29]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 149:40]
      host_lds_size_total_i <= 13'h0; // @[inflight_wg_buffer.scala 149:40]
    end else begin
      host_lds_size_total_i <= io_host_lds_size_total; // @[inflight_wg_buffer.scala 150:27]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 151:40]
      host_gds_size_total_i <= 11'h0; // @[inflight_wg_buffer.scala 151:40]
    end else begin
      host_gds_size_total_i <= io_host_gds_size_total; // @[inflight_wg_buffer.scala 152:27]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 153:47]
      dis_controller_start_alloc_i <= 1'h0; // @[inflight_wg_buffer.scala 153:47]
    end else begin
      dis_controller_start_alloc_i <= io_dis_controller_start_alloc; // @[inflight_wg_buffer.scala 154:34]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 155:50]
      dis_controller_wg_alloc_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 155:50]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      dis_controller_wg_alloc_valid_i <= _GEN_0;
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_wg_alloc_valid_i) begin // @[inflight_wg_buffer.scala 330:46]
        dis_controller_wg_alloc_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 331:43]
      end else begin
        dis_controller_wg_alloc_valid_i <= _GEN_0;
      end
    end else begin
      dis_controller_wg_alloc_valid_i <= _GEN_0;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 156:52]
      dis_controller_wg_dealloc_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 156:52]
    end else begin
      dis_controller_wg_dealloc_valid_i <= io_dis_controller_wg_dealloc_valid; // @[inflight_wg_buffer.scala 159:39]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 157:53]
      dis_controller_wg_rejected_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 157:53]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      dis_controller_wg_rejected_valid_i <= _GEN_2;
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_wg_alloc_valid_i) begin // @[inflight_wg_buffer.scala 330:46]
        dis_controller_wg_rejected_valid_i <= _GEN_2;
      end else begin
        dis_controller_wg_rejected_valid_i <= _GEN_36;
      end
    end else begin
      dis_controller_wg_rejected_valid_i <= _GEN_2;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 160:48]
      gpu_interface_dealloc_wg_id_i <= 5'h0; // @[inflight_wg_buffer.scala 160:48]
    end else begin
      gpu_interface_dealloc_wg_id_i <= io_gpu_interface_dealloc_wg_id; // @[inflight_wg_buffer.scala 161:35]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 162:40]
      inflight_tbl_alloc_st <= 8'h1; // @[inflight_wg_buffer.scala 162:40]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_start_alloc_i) begin // @[inflight_wg_buffer.scala 312:43]
        inflight_tbl_alloc_st <= 8'h2; // @[inflight_wg_buffer.scala 315:33]
      end else if (~wg_waiting_alloc_valid & (valid_not_pending_0 | valid_not_pending_1)) begin // @[inflight_wg_buffer.scala 317:81]
        inflight_tbl_alloc_st <= 8'h40; // @[inflight_wg_buffer.scala 318:33]
      end
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_wg_alloc_valid_i) begin // @[inflight_wg_buffer.scala 330:46]
        inflight_tbl_alloc_st <= 8'h4; // @[inflight_wg_buffer.scala 337:33]
      end else begin
        inflight_tbl_alloc_st <= _GEN_40;
      end
    end else if (8'h4 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      inflight_tbl_alloc_st <= _GEN_52;
    end else begin
      inflight_tbl_alloc_st <= _GEN_133;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 163:42]
      inflight_tbl_rd_host_st <= 4'h1; // @[inflight_wg_buffer.scala 163:42]
    end else if (4'h1 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
      if (host_wg_valid_i) begin // @[inflight_wg_buffer.scala 211:30]
        if (~waiting_tbl_valid_0 | ~waiting_tbl_valid_1) begin // @[inflight_wg_buffer.scala 212:52]
          inflight_tbl_rd_host_st <= 4'h2; // @[inflight_wg_buffer.scala 213:37]
        end
      end
    end else if (4'h2 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
      inflight_tbl_rd_host_st <= 4'h4; // @[inflight_wg_buffer.scala 225:33]
    end else if (4'h4 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
      inflight_tbl_rd_host_st <= 4'h8; // @[inflight_wg_buffer.scala 234:33]
    end else begin
      inflight_tbl_rd_host_st <= _GEN_10;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 164:40]
      allocator_wg_id_out_i <= 5'h0; // @[inflight_wg_buffer.scala 164:40]
    end else if (io_dis_controller_wg_rejected_valid) begin // @[inflight_wg_buffer.scala 169:46]
      allocator_wg_id_out_i <= io_allocator_wg_id_out; // @[inflight_wg_buffer.scala 171:29]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[inflight_wg_buffer.scala 165:43]
      allocator_wg_id_out_i <= io_allocator_wg_id_out; // @[inflight_wg_buffer.scala 167:29]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 173:52]
      inflight_wg_buffer_host_wf_done_i <= 1'h0; // @[inflight_wg_buffer.scala 173:52]
    end else begin
      inflight_wg_buffer_host_wf_done_i <= dis_controller_wg_dealloc_valid_i;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 175:58]
      inflight_wg_buffer_host_wf_done_wg_id_i <= 5'h0; // @[inflight_wg_buffer.scala 175:58]
    end else if (dis_controller_wg_dealloc_valid_i) begin // @[inflight_wg_buffer.scala 179:44]
      inflight_wg_buffer_host_wf_done_wg_id_i <= gpu_interface_dealloc_wg_id_i; // @[inflight_wg_buffer.scala 181:47]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 185:36]
      waiting_tbl_valid_0 <= 1'h0; // @[inflight_wg_buffer.scala 185:36]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      waiting_tbl_valid_0 <= _GEN_24;
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      waiting_tbl_valid_0 <= _GEN_24;
    end else if (8'h4 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      waiting_tbl_valid_0 <= _GEN_24;
    end else begin
      waiting_tbl_valid_0 <= _GEN_124;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 185:36]
      waiting_tbl_valid_1 <= 1'h0; // @[inflight_wg_buffer.scala 185:36]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      waiting_tbl_valid_1 <= _GEN_25;
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      waiting_tbl_valid_1 <= _GEN_25;
    end else if (8'h4 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      waiting_tbl_valid_1 <= _GEN_25;
    end else begin
      waiting_tbl_valid_1 <= _GEN_125;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 186:34]
      new_index_wr_en <= 1'h0; // @[inflight_wg_buffer.scala 186:34]
    end else if (4'h1 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
      new_index_wr_en <= 1'h0; // @[inflight_wg_buffer.scala 201:21]
    end else begin
      new_index_wr_en <= 4'h2 == inflight_tbl_rd_host_st;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 189:35]
      new_entry_wg_reg <= 58'h0; // @[inflight_wg_buffer.scala 189:35]
    end else if (!(4'h1 == inflight_tbl_rd_host_st)) begin // @[inflight_wg_buffer.scala 205:36]
      if (4'h2 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
        new_entry_wg_reg <= _new_entry_wg_reg_T; // @[inflight_wg_buffer.scala 223:26]
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 191:35]
      ready_tbl_wr_reg <= 73'h0; // @[inflight_wg_buffer.scala 191:35]
    end else if (!(4'h1 == inflight_tbl_rd_host_st)) begin // @[inflight_wg_buffer.scala 205:36]
      if (4'h2 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
        ready_tbl_wr_reg <= _ready_tbl_wr_reg_T; // @[inflight_wg_buffer.scala 224:26]
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 193:53]
      inflight_wg_buffer_host_rcvd_ack_i <= 1'h0; // @[inflight_wg_buffer.scala 193:53]
    end else if (4'h1 == inflight_tbl_rd_host_st) begin // @[inflight_wg_buffer.scala 205:36]
      inflight_wg_buffer_host_rcvd_ack_i <= 1'h0; // @[inflight_wg_buffer.scala 201:21]
    end else begin
      inflight_wg_buffer_host_rcvd_ack_i <= 4'h2 == inflight_tbl_rd_host_st;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 195:28]
      new_index <= 1'h0; // @[inflight_wg_buffer.scala 195:28]
    end else if (_T_1) begin // @[inflight_wg_buffer.scala 436:34]
      new_index <= 1'h0; // @[inflight_wg_buffer.scala 438:25]
    end else begin
      new_index <= _T_2;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 245:38]
      waiting_tbl_pending_0 <= 1'h0; // @[inflight_wg_buffer.scala 245:38]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_start_alloc_i) begin // @[inflight_wg_buffer.scala 312:43]
        waiting_tbl_pending_0 <= _GEN_27;
      end
    end else if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        waiting_tbl_pending_0 <= _GEN_126;
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 245:38]
      waiting_tbl_pending_1 <= 1'h0; // @[inflight_wg_buffer.scala 245:38]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_start_alloc_i) begin // @[inflight_wg_buffer.scala 312:43]
        waiting_tbl_pending_1 <= _GEN_28;
      end
    end else if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        waiting_tbl_pending_1 <= _GEN_127;
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 246:31]
      chosen_entry <= 1'h0; // @[inflight_wg_buffer.scala 246:31]
    end else if (waiting_tbl_valid_rotated_0) begin // @[inflight_wg_buffer.scala 460:41]
      chosen_entry <= _idx_found_entry_c_T_4[0] + 1'h1; // @[inflight_wg_buffer.scala 462:27]
    end else begin
      chosen_entry <= _GEN_226;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 247:44]
      chosen_entry_by_allocator <= 1'h0; // @[inflight_wg_buffer.scala 247:44]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          chosen_entry_by_allocator <= _GEN_136;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 248:40]
      chosen_entry_is_valid <= 1'h0; // @[inflight_wg_buffer.scala 248:40]
    end else begin
      chosen_entry_is_valid <= found_entry_valid_c; // @[inflight_wg_buffer.scala 430:27]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 249:32]
      wait_tbl_busy <= 1'h0; // @[inflight_wg_buffer.scala 249:32]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      wait_tbl_busy <= _GEN_35;
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      wait_tbl_busy <= 1'h0; // @[inflight_wg_buffer.scala 329:23]
    end else begin
      wait_tbl_busy <= 1'h1; // @[inflight_wg_buffer.scala 250:19]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 257:42]
      tbl_walk_wg_id_searched <= 5'h0; // @[inflight_wg_buffer.scala 257:42]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
        if (dis_controller_wg_alloc_valid_i) begin // @[inflight_wg_buffer.scala 330:46]
          tbl_walk_wg_id_searched <= allocator_wg_id_out_i; // @[inflight_wg_buffer.scala 332:35]
        end else begin
          tbl_walk_wg_id_searched <= _GEN_37;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 262:33]
      tbl_walk_rd_en <= 1'h0; // @[inflight_wg_buffer.scala 262:33]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      tbl_walk_rd_en <= 1'h0; // @[inflight_wg_buffer.scala 271:20]
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      tbl_walk_rd_en <= _GEN_43;
    end else if (8'h4 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      tbl_walk_rd_en <= _GEN_54;
    end else begin
      tbl_walk_rd_en <= _GEN_135;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 265:31]
      tbl_walk_idx <= 1'h0; // @[inflight_wg_buffer.scala 265:31]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
        if (dis_controller_wg_alloc_valid_i) begin // @[inflight_wg_buffer.scala 330:46]
          tbl_walk_idx <= 1'h0; // @[inflight_wg_buffer.scala 336:24]
        end else begin
          tbl_walk_idx <= _GEN_39;
        end
      end else if (8'h4 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
        tbl_walk_idx <= _GEN_53;
      end else begin
        tbl_walk_idx <= _GEN_134;
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 268:36]
      tbl_walk_rd_valid <= 1'h0; // @[inflight_wg_buffer.scala 268:36]
    end else begin
      tbl_walk_rd_valid <= tbl_walk_rd_en; // @[inflight_wg_buffer.scala 269:23]
    end
    if (reset) begin // @[inflight_wg_buffer.scala 274:49]
      inflight_wg_buffer_gpu_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 274:49]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      inflight_wg_buffer_gpu_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 305:36]
    end else if (8'h2 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      inflight_wg_buffer_gpu_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 305:36]
    end else if (8'h4 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      inflight_wg_buffer_gpu_valid_i <= 1'h0; // @[inflight_wg_buffer.scala 305:36]
    end else begin
      inflight_wg_buffer_gpu_valid_i <= 8'h8 == inflight_tbl_alloc_st;
    end
    if (reset) begin // @[inflight_wg_buffer.scala 276:60]
      inflight_wg_buffer_gpu_vgpr_size_per_wf_i <= 13'h0; // @[inflight_wg_buffer.scala 276:60]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_gpu_vgpr_size_per_wf_i <= _GEN_129;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 278:60]
      inflight_wg_buffer_gpu_sgpr_size_per_wf_i <= 13'h0; // @[inflight_wg_buffer.scala 278:60]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_gpu_sgpr_size_per_wf_i <= _GEN_130;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 280:51]
      inflight_wg_buffer_gpu_wf_size_i <= 10'h0; // @[inflight_wg_buffer.scala 280:51]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_gpu_wf_size_i <= _GEN_131;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 282:48]
      inflight_wg_buffer_start_pc_i <= 32'h0; // @[inflight_wg_buffer.scala 282:48]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_start_pc_i <= _GEN_132;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 286:51]
      inflight_wg_buffer_alloc_wg_id_i <= 5'h0; // @[inflight_wg_buffer.scala 286:51]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_alloc_wg_id_i <= _GEN_138;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 288:52]
      inflight_wg_buffer_alloc_num_wf_i <= 3'h0; // @[inflight_wg_buffer.scala 288:52]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_alloc_num_wf_i <= _GEN_139;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 290:55]
      inflight_wg_buffer_alloc_vgpr_size_i <= 13'h0; // @[inflight_wg_buffer.scala 290:55]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_alloc_vgpr_size_i <= _GEN_140;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 292:55]
      inflight_wg_buffer_alloc_sgpr_size_i <= 13'h0; // @[inflight_wg_buffer.scala 292:55]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_alloc_sgpr_size_i <= _GEN_141;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 294:54]
      inflight_wg_buffer_alloc_lds_size_i <= 13'h0; // @[inflight_wg_buffer.scala 294:54]
    end else if (!(8'h1 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
          inflight_wg_buffer_alloc_lds_size_i <= _GEN_142;
        end
      end
    end
    if (reset) begin // @[inflight_wg_buffer.scala 298:41]
      wg_waiting_alloc_valid <= 1'h0; // @[inflight_wg_buffer.scala 298:41]
    end else if (8'h1 == inflight_tbl_alloc_st) begin // @[inflight_wg_buffer.scala 306:34]
      if (dis_controller_start_alloc_i) begin // @[inflight_wg_buffer.scala 312:43]
        wg_waiting_alloc_valid <= 1'h0; // @[inflight_wg_buffer.scala 314:34]
      end
    end else if (!(8'h2 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
      if (!(8'h4 == inflight_tbl_alloc_st)) begin // @[inflight_wg_buffer.scala 306:34]
        wg_waiting_alloc_valid <= _GEN_137;
      end
    end
    last_chosen_entry_rr <= reset | _GEN_26; // @[inflight_wg_buffer.scala 300:{39,39}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  host_wg_valid_i = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  host_wg_id_i = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  host_num_wf_i = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  host_wf_size_i = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  host_start_pc_i = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  host_vgpr_size_total_i = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  host_sgpr_size_total_i = _RAND_6[12:0];
  _RAND_7 = {1{`RANDOM}};
  host_vgpr_size_per_wf_i = _RAND_7[12:0];
  _RAND_8 = {1{`RANDOM}};
  host_sgpr_size_per_wf_i = _RAND_8[12:0];
  _RAND_9 = {1{`RANDOM}};
  host_lds_size_total_i = _RAND_9[12:0];
  _RAND_10 = {1{`RANDOM}};
  host_gds_size_total_i = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  dis_controller_start_alloc_i = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dis_controller_wg_alloc_valid_i = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  dis_controller_wg_dealloc_valid_i = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dis_controller_wg_rejected_valid_i = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  gpu_interface_dealloc_wg_id_i = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  inflight_tbl_alloc_st = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_tbl_rd_host_st = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  allocator_wg_id_out_i = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_wg_buffer_host_wf_done_i = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inflight_wg_buffer_host_wf_done_wg_id_i = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  waiting_tbl_valid_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  waiting_tbl_valid_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  new_index_wr_en = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  new_entry_wg_reg = _RAND_24[57:0];
  _RAND_25 = {3{`RANDOM}};
  ready_tbl_wr_reg = _RAND_25[72:0];
  _RAND_26 = {1{`RANDOM}};
  inflight_wg_buffer_host_rcvd_ack_i = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  new_index = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  waiting_tbl_pending_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  waiting_tbl_pending_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  chosen_entry = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  chosen_entry_by_allocator = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  chosen_entry_is_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  wait_tbl_busy = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tbl_walk_wg_id_searched = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  tbl_walk_rd_en = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tbl_walk_idx = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  tbl_walk_rd_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_valid_i = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_vgpr_size_per_wf_i = _RAND_39[12:0];
  _RAND_40 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_sgpr_size_per_wf_i = _RAND_40[12:0];
  _RAND_41 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_wf_size_i = _RAND_41[9:0];
  _RAND_42 = {1{`RANDOM}};
  inflight_wg_buffer_start_pc_i = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  inflight_wg_buffer_alloc_wg_id_i = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  inflight_wg_buffer_alloc_num_wf_i = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  inflight_wg_buffer_alloc_vgpr_size_i = _RAND_45[12:0];
  _RAND_46 = {1{`RANDOM}};
  inflight_wg_buffer_alloc_sgpr_size_i = _RAND_46[12:0];
  _RAND_47 = {1{`RANDOM}};
  inflight_wg_buffer_alloc_lds_size_i = _RAND_47[12:0];
  _RAND_48 = {1{`RANDOM}};
  wg_waiting_alloc_valid = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  last_chosen_entry_rr = _RAND_49[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_2(
  input        clock,
  input        reset,
  input  [1:0] io_rd_addr,
  input  [1:0] io_wr_addr,
  input  [7:0] io_wr_word,
  output [7:0] io_rd_word,
  input        io_wr_en,
  input        io_rd_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:3]; // @[RAM.scala 14:18]
  wire  mem_rd_word_reg_MPORT_en; // @[RAM.scala 14:18]
  wire [1:0] mem_rd_word_reg_MPORT_addr; // @[RAM.scala 14:18]
  wire [7:0] mem_rd_word_reg_MPORT_data; // @[RAM.scala 14:18]
  wire [7:0] mem_MPORT_data; // @[RAM.scala 14:18]
  wire [1:0] mem_MPORT_addr; // @[RAM.scala 14:18]
  wire  mem_MPORT_mask; // @[RAM.scala 14:18]
  wire  mem_MPORT_en; // @[RAM.scala 14:18]
  reg [7:0] rd_word_reg; // @[RAM.scala 19:30]
  assign mem_rd_word_reg_MPORT_en = io_rd_en;
  assign mem_rd_word_reg_MPORT_addr = io_rd_addr;
  assign mem_rd_word_reg_MPORT_data = mem[mem_rd_word_reg_MPORT_addr]; // @[RAM.scala 14:18]
  assign mem_MPORT_data = io_wr_word;
  assign mem_MPORT_addr = io_wr_addr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wr_en;
  assign io_rd_word = rd_word_reg; // @[RAM.scala 23:16]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[RAM.scala 14:18]
    end
    if (reset) begin // @[RAM.scala 19:30]
      rd_word_reg <= 8'h0; // @[RAM.scala 19:30]
    end else if (io_rd_en) begin // @[RAM.scala 20:20]
      rd_word_reg <= mem_rd_word_reg_MPORT_data; // @[RAM.scala 21:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rd_word_reg = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cu_handler(
  input        clock,
  input        reset,
  input        io_wg_alloc_en,
  input  [4:0] io_wg_alloc_wg_id,
  input  [2:0] io_wg_alloc_wf_count,
  input        io_ready_for_dispatch2cu,
  output       io_dispatch2cu_wf_dispatch,
  output [4:0] io_dispatch2cu_wf_tag_dispatch,
  input        io_cu2dispatch_wf_done_i,
  input  [4:0] io_cu2dispatch_wf_tag_done_i,
  input        io_wg_done_ack,
  output       io_wg_done_valid,
  output [4:0] io_wg_done_wg_id,
  output       io_invalid_due_to_not_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  info_ram_clock; // @[cu_handler.scala 108:26]
  wire  info_ram_reset; // @[cu_handler.scala 108:26]
  wire [1:0] info_ram_io_rd_addr; // @[cu_handler.scala 108:26]
  wire [1:0] info_ram_io_wr_addr; // @[cu_handler.scala 108:26]
  wire [7:0] info_ram_io_wr_word; // @[cu_handler.scala 108:26]
  wire [7:0] info_ram_io_rd_word; // @[cu_handler.scala 108:26]
  wire  info_ram_io_wr_en; // @[cu_handler.scala 108:26]
  wire  info_ram_io_rd_en; // @[cu_handler.scala 108:26]
  reg [1:0] next_free_slot; // @[cu_handler.scala 35:33]
  reg  used_slot_bitmap_0; // @[cu_handler.scala 37:35]
  reg  used_slot_bitmap_1; // @[cu_handler.scala 37:35]
  reg  used_slot_bitmap_2; // @[cu_handler.scala 37:35]
  reg  used_slot_bitmap_3; // @[cu_handler.scala 37:35]
  reg  pending_wg_bitmap_0; // @[cu_handler.scala 38:36]
  reg  pending_wg_bitmap_1; // @[cu_handler.scala 38:36]
  reg  pending_wg_bitmap_2; // @[cu_handler.scala 38:36]
  reg  pending_wg_bitmap_3; // @[cu_handler.scala 38:36]
  reg [2:0] pending_wf_count_0; // @[cu_handler.scala 48:35]
  reg [2:0] pending_wf_count_1; // @[cu_handler.scala 48:35]
  reg [2:0] pending_wf_count_2; // @[cu_handler.scala 48:35]
  reg [2:0] pending_wf_count_3; // @[cu_handler.scala 48:35]
  reg [2:0] curr_alloc_wf_count; // @[cu_handler.scala 49:38]
  reg [1:0] curr_alloc_wf_slot; // @[cu_handler.scala 50:37]
  reg  dispatch2cu_wf_dispatch_i; // @[cu_handler.scala 51:44]
  reg [4:0] dispatch2cu_wf_tag_dispatch_i; // @[cu_handler.scala 52:48]
  reg  next_served_dealloc_valid; // @[cu_handler.scala 59:44]
  reg [1:0] next_served_dealloc; // @[cu_handler.scala 61:38]
  reg [1:0] curr_dealloc_wg_slot; // @[cu_handler.scala 71:39]
  reg  info_ram_rd_en; // @[cu_handler.scala 74:33]
  reg  info_ram_rd_valid; // @[cu_handler.scala 75:36]
  reg  info_ram_wr_en; // @[cu_handler.scala 77:33]
  reg [1:0] info_ram_wr_addr; // @[cu_handler.scala 78:35]
  reg [7:0] info_ram_wr_reg; // @[cu_handler.scala 79:34]
  reg  wg_done_valid_i; // @[cu_handler.scala 80:34]
  reg [4:0] wg_done_wg_id_i; // @[cu_handler.scala 81:34]
  reg [2:0] curr_wf_count; // @[cu_handler.scala 82:32]
  reg [1:0] alloc_st; // @[cu_handler.scala 87:27]
  reg [2:0] dealloc_st; // @[cu_handler.scala 93:29]
  reg  invalid_due_to_not_ready_i; // @[cu_handler.scala 116:45]
  reg  next_free_slot_valid; // @[cu_handler.scala 121:39]
  wire  _T_1 = io_wg_alloc_en & next_free_slot_valid; // @[cu_handler.scala 129:33]
  wire [7:0] _info_ram_wr_reg_T = {io_wg_alloc_wg_id,io_wg_alloc_wf_count}; // @[Cat.scala 31:58]
  wire  _GEN_0 = 2'h0 == next_free_slot | used_slot_bitmap_0; // @[cu_handler.scala 135:{50,50} 37:35]
  wire  _GEN_1 = 2'h1 == next_free_slot | used_slot_bitmap_1; // @[cu_handler.scala 135:{50,50} 37:35]
  wire  _GEN_2 = 2'h2 == next_free_slot | used_slot_bitmap_2; // @[cu_handler.scala 135:{50,50} 37:35]
  wire  _GEN_3 = 2'h3 == next_free_slot | used_slot_bitmap_3; // @[cu_handler.scala 135:{50,50} 37:35]
  wire [2:0] _GEN_4 = 2'h0 == next_free_slot ? io_wg_alloc_wf_count : pending_wf_count_0; // @[cu_handler.scala 137:{50,50} 48:35]
  wire [2:0] _GEN_5 = 2'h1 == next_free_slot ? io_wg_alloc_wf_count : pending_wf_count_1; // @[cu_handler.scala 137:{50,50} 48:35]
  wire [2:0] _GEN_6 = 2'h2 == next_free_slot ? io_wg_alloc_wf_count : pending_wf_count_2; // @[cu_handler.scala 137:{50,50} 48:35]
  wire [2:0] _GEN_7 = 2'h3 == next_free_slot ? io_wg_alloc_wf_count : pending_wf_count_3; // @[cu_handler.scala 137:{50,50} 48:35]
  wire  _GEN_13 = io_wg_alloc_en & next_free_slot_valid ? _GEN_0 : used_slot_bitmap_0; // @[cu_handler.scala 129:57 37:35]
  wire  _GEN_14 = io_wg_alloc_en & next_free_slot_valid ? _GEN_1 : used_slot_bitmap_1; // @[cu_handler.scala 129:57 37:35]
  wire  _GEN_15 = io_wg_alloc_en & next_free_slot_valid ? _GEN_2 : used_slot_bitmap_2; // @[cu_handler.scala 129:57 37:35]
  wire  _GEN_16 = io_wg_alloc_en & next_free_slot_valid ? _GEN_3 : used_slot_bitmap_3; // @[cu_handler.scala 129:57 37:35]
  wire [2:0] _GEN_17 = io_wg_alloc_en & next_free_slot_valid ? _GEN_4 : pending_wf_count_0; // @[cu_handler.scala 129:57 48:35]
  wire [2:0] _GEN_18 = io_wg_alloc_en & next_free_slot_valid ? _GEN_5 : pending_wf_count_1; // @[cu_handler.scala 129:57 48:35]
  wire [2:0] _GEN_19 = io_wg_alloc_en & next_free_slot_valid ? _GEN_6 : pending_wf_count_2; // @[cu_handler.scala 129:57 48:35]
  wire [2:0] _GEN_20 = io_wg_alloc_en & next_free_slot_valid ? _GEN_7 : pending_wf_count_3; // @[cu_handler.scala 129:57 48:35]
  wire [2:0] _dispatch2cu_wf_tag_dispatch_i_T_1 = curr_alloc_wf_count - 3'h1; // @[cu_handler.scala 147:98]
  wire [4:0] _dispatch2cu_wf_tag_dispatch_i_T_2 = {curr_alloc_wf_slot,_dispatch2cu_wf_tag_dispatch_i_T_1}; // @[Cat.scala 31:58]
  wire [4:0] _GEN_23 = io_ready_for_dispatch2cu ? _dispatch2cu_wf_tag_dispatch_i_T_2 : dispatch2cu_wf_tag_dispatch_i; // @[cu_handler.scala 143:47 147:51 52:48]
  wire [2:0] _GEN_24 = io_ready_for_dispatch2cu ? _dispatch2cu_wf_tag_dispatch_i_T_1 : curr_alloc_wf_count; // @[cu_handler.scala 143:47 148:41 49:38]
  wire  _GEN_25 = io_ready_for_dispatch2cu ? 1'h0 : 1'h1; // @[cu_handler.scala 143:47 149:48 153:48]
  wire  _GEN_26 = curr_alloc_wf_count != 3'h0 & io_ready_for_dispatch2cu; // @[cu_handler.scala 123:31 142:46]
  wire  _GEN_29 = curr_alloc_wf_count != 3'h0 & _GEN_25; // @[cu_handler.scala 142:46 158:44]
  wire  _GEN_36 = 2'h1 == alloc_st & _T_1; // @[cu_handler.scala 118:20 127:21]
  wire  _GEN_41 = 2'h1 == alloc_st ? _GEN_13 : used_slot_bitmap_0; // @[cu_handler.scala 127:21 37:35]
  wire  _GEN_42 = 2'h1 == alloc_st ? _GEN_14 : used_slot_bitmap_1; // @[cu_handler.scala 127:21 37:35]
  wire  _GEN_43 = 2'h1 == alloc_st ? _GEN_15 : used_slot_bitmap_2; // @[cu_handler.scala 127:21 37:35]
  wire  _GEN_44 = 2'h1 == alloc_st ? _GEN_16 : used_slot_bitmap_3; // @[cu_handler.scala 127:21 37:35]
  wire [2:0] _GEN_45 = 2'h1 == alloc_st ? _GEN_17 : pending_wf_count_0; // @[cu_handler.scala 127:21 48:35]
  wire [2:0] _GEN_46 = 2'h1 == alloc_st ? _GEN_18 : pending_wf_count_1; // @[cu_handler.scala 127:21 48:35]
  wire [2:0] _GEN_47 = 2'h1 == alloc_st ? _GEN_19 : pending_wf_count_2; // @[cu_handler.scala 127:21 48:35]
  wire [2:0] _GEN_48 = 2'h1 == alloc_st ? _GEN_20 : pending_wf_count_3; // @[cu_handler.scala 127:21 48:35]
  wire [2:0] _GEN_54 = 2'h1 == next_served_dealloc ? pending_wf_count_1 : pending_wf_count_0; // @[cu_handler.scala 174:{31,31}]
  wire [2:0] _GEN_55 = 2'h2 == next_served_dealloc ? pending_wf_count_2 : _GEN_54; // @[cu_handler.scala 174:{31,31}]
  wire  _GEN_57 = 2'h0 == next_served_dealloc ? 1'h0 : pending_wg_bitmap_0; // @[cu_handler.scala 175:{56,56} 38:36]
  wire  _GEN_58 = 2'h1 == next_served_dealloc ? 1'h0 : pending_wg_bitmap_1; // @[cu_handler.scala 175:{56,56} 38:36]
  wire  _GEN_59 = 2'h2 == next_served_dealloc ? 1'h0 : pending_wg_bitmap_2; // @[cu_handler.scala 175:{56,56} 38:36]
  wire  _GEN_60 = 2'h3 == next_served_dealloc ? 1'h0 : pending_wg_bitmap_3; // @[cu_handler.scala 175:{56,56} 38:36]
  wire  _GEN_64 = next_served_dealloc_valid ? _GEN_57 : pending_wg_bitmap_0; // @[cu_handler.scala 171:44 38:36]
  wire  _GEN_65 = next_served_dealloc_valid ? _GEN_58 : pending_wg_bitmap_1; // @[cu_handler.scala 171:44 38:36]
  wire  _GEN_66 = next_served_dealloc_valid ? _GEN_59 : pending_wg_bitmap_2; // @[cu_handler.scala 171:44 38:36]
  wire  _GEN_67 = next_served_dealloc_valid ? _GEN_60 : pending_wg_bitmap_3; // @[cu_handler.scala 171:44 38:36]
  wire  _T_6 = curr_wf_count == 3'h0; // @[cu_handler.scala 181:36]
  wire [7:0] info_ram_rd_reg = info_ram_io_rd_word; // @[cu_handler.scala 114:21 76:31]
  wire  _GEN_69 = 2'h0 == curr_dealloc_wg_slot ? 1'h0 : _GEN_41; // @[cu_handler.scala 184:{60,60}]
  wire  _GEN_70 = 2'h1 == curr_dealloc_wg_slot ? 1'h0 : _GEN_42; // @[cu_handler.scala 184:{60,60}]
  wire  _GEN_71 = 2'h2 == curr_dealloc_wg_slot ? 1'h0 : _GEN_43; // @[cu_handler.scala 184:{60,60}]
  wire  _GEN_72 = 2'h3 == curr_dealloc_wg_slot ? 1'h0 : _GEN_44; // @[cu_handler.scala 184:{60,60}]
  wire [4:0] _GEN_74 = curr_wf_count == 3'h0 ? info_ram_rd_reg[7:3] : wg_done_wg_id_i; // @[cu_handler.scala 181:44 183:37 81:34]
  wire  _GEN_75 = curr_wf_count == 3'h0 ? _GEN_69 : _GEN_41; // @[cu_handler.scala 181:44]
  wire  _GEN_76 = curr_wf_count == 3'h0 ? _GEN_70 : _GEN_42; // @[cu_handler.scala 181:44]
  wire  _GEN_77 = curr_wf_count == 3'h0 ? _GEN_71 : _GEN_43; // @[cu_handler.scala 181:44]
  wire  _GEN_78 = curr_wf_count == 3'h0 ? _GEN_72 : _GEN_44; // @[cu_handler.scala 181:44]
  wire [2:0] _GEN_79 = curr_wf_count == 3'h0 ? 3'h4 : 3'h1; // @[cu_handler.scala 181:44 185:32 188:32]
  wire  _GEN_80 = info_ram_rd_valid & _T_6; // @[cu_handler.scala 166:21 180:36]
  wire [2:0] _GEN_87 = io_wg_done_ack ? 3'h1 : dealloc_st; // @[cu_handler.scala 193:33 194:28 93:29]
  wire  _GEN_88 = io_wg_done_ack ? 1'h0 : 1'h1; // @[cu_handler.scala 166:21 193:33 197:33]
  wire  _GEN_90 = 3'h4 == dealloc_st & _GEN_88; // @[cu_handler.scala 166:21 169:23]
  wire  _GEN_98 = 3'h1 == dealloc_st & next_served_dealloc_valid; // @[cu_handler.scala 164:20 169:23]
  wire  _GEN_101 = 3'h1 == dealloc_st ? _GEN_64 : pending_wg_bitmap_0; // @[cu_handler.scala 169:23 38:36]
  wire  _GEN_102 = 3'h1 == dealloc_st ? _GEN_65 : pending_wg_bitmap_1; // @[cu_handler.scala 169:23 38:36]
  wire  _GEN_103 = 3'h1 == dealloc_st ? _GEN_66 : pending_wg_bitmap_2; // @[cu_handler.scala 169:23 38:36]
  wire  _GEN_104 = 3'h1 == dealloc_st ? _GEN_67 : pending_wg_bitmap_3; // @[cu_handler.scala 169:23 38:36]
  wire  _GEN_112 = 2'h0 == io_cu2dispatch_wf_tag_done_i[4:3] | _GEN_101; // @[cu_handler.scala 202:{93,93}]
  wire  _GEN_113 = 2'h1 == io_cu2dispatch_wf_tag_done_i[4:3] | _GEN_102; // @[cu_handler.scala 202:{93,93}]
  wire  _GEN_114 = 2'h2 == io_cu2dispatch_wf_tag_done_i[4:3] | _GEN_103; // @[cu_handler.scala 202:{93,93}]
  wire  _GEN_115 = 2'h3 == io_cu2dispatch_wf_tag_done_i[4:3] | _GEN_104; // @[cu_handler.scala 202:{93,93}]
  wire [2:0] _GEN_117 = 2'h1 == io_cu2dispatch_wf_tag_done_i[4:3] ? pending_wf_count_1 : pending_wf_count_0; // @[cu_handler.scala 204:{178,178}]
  wire [2:0] _GEN_118 = 2'h2 == io_cu2dispatch_wf_tag_done_i[4:3] ? pending_wf_count_2 : _GEN_117; // @[cu_handler.scala 204:{178,178}]
  wire [2:0] _GEN_119 = 2'h3 == io_cu2dispatch_wf_tag_done_i[4:3] ? pending_wf_count_3 : _GEN_118; // @[cu_handler.scala 204:{178,178}]
  wire [2:0] _pending_wf_count_T_2 = _GEN_119 - 3'h1; // @[cu_handler.scala 204:178]
  wire [1:0] _GEN_133 = pending_wg_bitmap_3 ? 2'h3 : 2'h0; // @[cu_handler.scala 216:24 218:35 220:32]
  wire  found_free_slot_valid = pending_wg_bitmap_0 | (pending_wg_bitmap_1 | (pending_wg_bitmap_2 | pending_wg_bitmap_3)
    ); // @[cu_handler.scala 218:35 219:35]
  wire [1:0] _GEN_141 = ~used_slot_bitmap_3 ? 2'h3 : 2'h0; // @[cu_handler.scala 230:25 232:35 234:33]
  wire  found_free_slot_valid2 = ~used_slot_bitmap_0 | (~used_slot_bitmap_1 | (~used_slot_bitmap_2 | ~used_slot_bitmap_3
    )); // @[cu_handler.scala 232:35 233:36]
  RAM_2 info_ram ( // @[cu_handler.scala 108:26]
    .clock(info_ram_clock),
    .reset(info_ram_reset),
    .io_rd_addr(info_ram_io_rd_addr),
    .io_wr_addr(info_ram_io_wr_addr),
    .io_wr_word(info_ram_io_wr_word),
    .io_rd_word(info_ram_io_rd_word),
    .io_wr_en(info_ram_io_wr_en),
    .io_rd_en(info_ram_io_rd_en)
  );
  assign io_dispatch2cu_wf_dispatch = dispatch2cu_wf_dispatch_i; // @[cu_handler.scala 206:32]
  assign io_dispatch2cu_wf_tag_dispatch = dispatch2cu_wf_tag_dispatch_i; // @[cu_handler.scala 207:36]
  assign io_wg_done_valid = wg_done_valid_i; // @[cu_handler.scala 209:22]
  assign io_wg_done_wg_id = wg_done_wg_id_i; // @[cu_handler.scala 210:22]
  assign io_invalid_due_to_not_ready = invalid_due_to_not_ready_i; // @[cu_handler.scala 238:33]
  assign info_ram_clock = clock;
  assign info_ram_reset = reset;
  assign info_ram_io_rd_addr = curr_dealloc_wg_slot; // @[cu_handler.scala 113:25]
  assign info_ram_io_wr_addr = info_ram_wr_addr; // @[cu_handler.scala 110:25]
  assign info_ram_io_wr_word = info_ram_wr_reg; // @[cu_handler.scala 111:25]
  assign info_ram_io_wr_en = info_ram_wr_en; // @[cu_handler.scala 109:23]
  assign info_ram_io_rd_en = info_ram_rd_en; // @[cu_handler.scala 112:23]
  always @(posedge clock) begin
    if (reset) begin // @[cu_handler.scala 35:33]
      next_free_slot <= 2'h0; // @[cu_handler.scala 35:33]
    end else if (~used_slot_bitmap_0) begin // @[cu_handler.scala 232:35]
      next_free_slot <= 2'h0; // @[cu_handler.scala 234:33]
    end else if (~used_slot_bitmap_1) begin // @[cu_handler.scala 232:35]
      next_free_slot <= 2'h1; // @[cu_handler.scala 234:33]
    end else if (~used_slot_bitmap_2) begin // @[cu_handler.scala 232:35]
      next_free_slot <= 2'h2; // @[cu_handler.scala 234:33]
    end else begin
      next_free_slot <= _GEN_141;
    end
    if (reset) begin // @[cu_handler.scala 37:35]
      used_slot_bitmap_0 <= 1'h0; // @[cu_handler.scala 37:35]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      used_slot_bitmap_0 <= _GEN_41;
    end else if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (info_ram_rd_valid) begin // @[cu_handler.scala 180:36]
        used_slot_bitmap_0 <= _GEN_75;
      end else begin
        used_slot_bitmap_0 <= _GEN_41;
      end
    end else begin
      used_slot_bitmap_0 <= _GEN_41;
    end
    if (reset) begin // @[cu_handler.scala 37:35]
      used_slot_bitmap_1 <= 1'h0; // @[cu_handler.scala 37:35]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      used_slot_bitmap_1 <= _GEN_42;
    end else if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (info_ram_rd_valid) begin // @[cu_handler.scala 180:36]
        used_slot_bitmap_1 <= _GEN_76;
      end else begin
        used_slot_bitmap_1 <= _GEN_42;
      end
    end else begin
      used_slot_bitmap_1 <= _GEN_42;
    end
    if (reset) begin // @[cu_handler.scala 37:35]
      used_slot_bitmap_2 <= 1'h0; // @[cu_handler.scala 37:35]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      used_slot_bitmap_2 <= _GEN_43;
    end else if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (info_ram_rd_valid) begin // @[cu_handler.scala 180:36]
        used_slot_bitmap_2 <= _GEN_77;
      end else begin
        used_slot_bitmap_2 <= _GEN_43;
      end
    end else begin
      used_slot_bitmap_2 <= _GEN_43;
    end
    if (reset) begin // @[cu_handler.scala 37:35]
      used_slot_bitmap_3 <= 1'h0; // @[cu_handler.scala 37:35]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      used_slot_bitmap_3 <= _GEN_44;
    end else if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (info_ram_rd_valid) begin // @[cu_handler.scala 180:36]
        used_slot_bitmap_3 <= _GEN_78;
      end else begin
        used_slot_bitmap_3 <= _GEN_44;
      end
    end else begin
      used_slot_bitmap_3 <= _GEN_44;
    end
    if (reset) begin // @[cu_handler.scala 38:36]
      pending_wg_bitmap_0 <= 1'h0; // @[cu_handler.scala 38:36]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      pending_wg_bitmap_0 <= _GEN_112;
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        pending_wg_bitmap_0 <= _GEN_57;
      end
    end
    if (reset) begin // @[cu_handler.scala 38:36]
      pending_wg_bitmap_1 <= 1'h0; // @[cu_handler.scala 38:36]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      pending_wg_bitmap_1 <= _GEN_113;
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        pending_wg_bitmap_1 <= _GEN_58;
      end
    end
    if (reset) begin // @[cu_handler.scala 38:36]
      pending_wg_bitmap_2 <= 1'h0; // @[cu_handler.scala 38:36]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      pending_wg_bitmap_2 <= _GEN_114;
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        pending_wg_bitmap_2 <= _GEN_59;
      end
    end
    if (reset) begin // @[cu_handler.scala 38:36]
      pending_wg_bitmap_3 <= 1'h0; // @[cu_handler.scala 38:36]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      pending_wg_bitmap_3 <= _GEN_115;
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        pending_wg_bitmap_3 <= _GEN_60;
      end
    end
    if (reset) begin // @[cu_handler.scala 48:35]
      pending_wf_count_0 <= 3'h0; // @[cu_handler.scala 48:35]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      if (2'h0 == io_cu2dispatch_wf_tag_done_i[4:3]) begin // @[cu_handler.scala 204:92]
        pending_wf_count_0 <= _pending_wf_count_T_2; // @[cu_handler.scala 204:92]
      end else begin
        pending_wf_count_0 <= _GEN_45;
      end
    end else begin
      pending_wf_count_0 <= _GEN_45;
    end
    if (reset) begin // @[cu_handler.scala 48:35]
      pending_wf_count_1 <= 3'h0; // @[cu_handler.scala 48:35]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      if (2'h1 == io_cu2dispatch_wf_tag_done_i[4:3]) begin // @[cu_handler.scala 204:92]
        pending_wf_count_1 <= _pending_wf_count_T_2; // @[cu_handler.scala 204:92]
      end else begin
        pending_wf_count_1 <= _GEN_46;
      end
    end else begin
      pending_wf_count_1 <= _GEN_46;
    end
    if (reset) begin // @[cu_handler.scala 48:35]
      pending_wf_count_2 <= 3'h0; // @[cu_handler.scala 48:35]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      if (2'h2 == io_cu2dispatch_wf_tag_done_i[4:3]) begin // @[cu_handler.scala 204:92]
        pending_wf_count_2 <= _pending_wf_count_T_2; // @[cu_handler.scala 204:92]
      end else begin
        pending_wf_count_2 <= _GEN_47;
      end
    end else begin
      pending_wf_count_2 <= _GEN_47;
    end
    if (reset) begin // @[cu_handler.scala 48:35]
      pending_wf_count_3 <= 3'h0; // @[cu_handler.scala 48:35]
    end else if (io_cu2dispatch_wf_done_i) begin // @[cu_handler.scala 201:35]
      if (2'h3 == io_cu2dispatch_wf_tag_done_i[4:3]) begin // @[cu_handler.scala 204:92]
        pending_wf_count_3 <= _pending_wf_count_T_2; // @[cu_handler.scala 204:92]
      end else begin
        pending_wf_count_3 <= _GEN_48;
      end
    end else begin
      pending_wf_count_3 <= _GEN_48;
    end
    if (reset) begin // @[cu_handler.scala 49:38]
      curr_alloc_wf_count <= 3'h0; // @[cu_handler.scala 49:38]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (io_wg_alloc_en & next_free_slot_valid) begin // @[cu_handler.scala 129:57]
        curr_alloc_wf_count <= io_wg_alloc_wf_count; // @[cu_handler.scala 133:37]
      end
    end else if (2'h2 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (curr_alloc_wf_count != 3'h0) begin // @[cu_handler.scala 142:46]
        curr_alloc_wf_count <= _GEN_24;
      end
    end
    if (reset) begin // @[cu_handler.scala 50:37]
      curr_alloc_wf_slot <= 2'h0; // @[cu_handler.scala 50:37]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (io_wg_alloc_en & next_free_slot_valid) begin // @[cu_handler.scala 129:57]
        curr_alloc_wf_slot <= next_free_slot; // @[cu_handler.scala 134:36]
      end
    end
    if (reset) begin // @[cu_handler.scala 51:44]
      dispatch2cu_wf_dispatch_i <= 1'h0; // @[cu_handler.scala 51:44]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      dispatch2cu_wf_dispatch_i <= 1'h0; // @[cu_handler.scala 123:31]
    end else begin
      dispatch2cu_wf_dispatch_i <= 2'h2 == alloc_st & _GEN_26;
    end
    if (reset) begin // @[cu_handler.scala 52:48]
      dispatch2cu_wf_tag_dispatch_i <= 5'h0; // @[cu_handler.scala 52:48]
    end else if (!(2'h1 == alloc_st)) begin // @[cu_handler.scala 127:21]
      if (2'h2 == alloc_st) begin // @[cu_handler.scala 127:21]
        if (curr_alloc_wf_count != 3'h0) begin // @[cu_handler.scala 142:46]
          dispatch2cu_wf_tag_dispatch_i <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[cu_handler.scala 59:44]
      next_served_dealloc_valid <= 1'h0; // @[cu_handler.scala 59:44]
    end else begin
      next_served_dealloc_valid <= found_free_slot_valid; // @[cu_handler.scala 162:31]
    end
    if (reset) begin // @[cu_handler.scala 61:38]
      next_served_dealloc <= 2'h0; // @[cu_handler.scala 61:38]
    end else if (pending_wg_bitmap_0) begin // @[cu_handler.scala 218:35]
      next_served_dealloc <= 2'h0; // @[cu_handler.scala 220:32]
    end else if (pending_wg_bitmap_1) begin // @[cu_handler.scala 218:35]
      next_served_dealloc <= 2'h1; // @[cu_handler.scala 220:32]
    end else if (pending_wg_bitmap_2) begin // @[cu_handler.scala 218:35]
      next_served_dealloc <= 2'h2; // @[cu_handler.scala 220:32]
    end else begin
      next_served_dealloc <= _GEN_133;
    end
    if (reset) begin // @[cu_handler.scala 71:39]
      curr_dealloc_wg_slot <= 2'h0; // @[cu_handler.scala 71:39]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        curr_dealloc_wg_slot <= next_served_dealloc; // @[cu_handler.scala 173:38]
      end
    end
    if (reset) begin // @[cu_handler.scala 74:33]
      info_ram_rd_en <= 1'h0; // @[cu_handler.scala 74:33]
    end else begin
      info_ram_rd_en <= _GEN_98;
    end
    if (reset) begin // @[cu_handler.scala 75:36]
      info_ram_rd_valid <= 1'h0; // @[cu_handler.scala 75:36]
    end else begin
      info_ram_rd_valid <= info_ram_rd_en; // @[cu_handler.scala 165:23]
    end
    if (reset) begin // @[cu_handler.scala 77:33]
      info_ram_wr_en <= 1'h0; // @[cu_handler.scala 77:33]
    end else begin
      info_ram_wr_en <= _GEN_36;
    end
    if (reset) begin // @[cu_handler.scala 78:35]
      info_ram_wr_addr <= 2'h0; // @[cu_handler.scala 78:35]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (io_wg_alloc_en & next_free_slot_valid) begin // @[cu_handler.scala 129:57]
        info_ram_wr_addr <= next_free_slot; // @[cu_handler.scala 131:34]
      end
    end
    if (reset) begin // @[cu_handler.scala 79:34]
      info_ram_wr_reg <= 8'h0; // @[cu_handler.scala 79:34]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (io_wg_alloc_en & next_free_slot_valid) begin // @[cu_handler.scala 129:57]
        info_ram_wr_reg <= _info_ram_wr_reg_T; // @[cu_handler.scala 132:33]
      end
    end
    if (reset) begin // @[cu_handler.scala 80:34]
      wg_done_valid_i <= 1'h0; // @[cu_handler.scala 80:34]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      wg_done_valid_i <= 1'h0; // @[cu_handler.scala 166:21]
    end else if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
      wg_done_valid_i <= _GEN_80;
    end else begin
      wg_done_valid_i <= _GEN_90;
    end
    if (reset) begin // @[cu_handler.scala 81:34]
      wg_done_wg_id_i <= 5'h0; // @[cu_handler.scala 81:34]
    end else if (!(3'h1 == dealloc_st)) begin // @[cu_handler.scala 169:23]
      if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
        if (info_ram_rd_valid) begin // @[cu_handler.scala 180:36]
          wg_done_wg_id_i <= _GEN_74;
        end
      end
    end
    if (reset) begin // @[cu_handler.scala 82:32]
      curr_wf_count <= 3'h0; // @[cu_handler.scala 82:32]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        if (2'h3 == next_served_dealloc) begin // @[cu_handler.scala 174:31]
          curr_wf_count <= pending_wf_count_3; // @[cu_handler.scala 174:31]
        end else begin
          curr_wf_count <= _GEN_55;
        end
      end
    end
    if (reset) begin // @[cu_handler.scala 87:27]
      alloc_st <= 2'h1; // @[cu_handler.scala 87:27]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (io_wg_alloc_en & next_free_slot_valid) begin // @[cu_handler.scala 129:57]
        alloc_st <= 2'h2; // @[cu_handler.scala 138:26]
      end
    end else if (2'h2 == alloc_st) begin // @[cu_handler.scala 127:21]
      if (!(curr_alloc_wf_count != 3'h0)) begin // @[cu_handler.scala 142:46]
        alloc_st <= 2'h1; // @[cu_handler.scala 157:26]
      end
    end
    if (reset) begin // @[cu_handler.scala 93:29]
      dealloc_st <= 3'h1; // @[cu_handler.scala 93:29]
    end else if (3'h1 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (next_served_dealloc_valid) begin // @[cu_handler.scala 171:44]
        dealloc_st <= 3'h2; // @[cu_handler.scala 176:28]
      end
    end else if (3'h2 == dealloc_st) begin // @[cu_handler.scala 169:23]
      if (info_ram_rd_valid) begin // @[cu_handler.scala 180:36]
        dealloc_st <= _GEN_79;
      end
    end else if (3'h4 == dealloc_st) begin // @[cu_handler.scala 169:23]
      dealloc_st <= _GEN_87;
    end
    if (reset) begin // @[cu_handler.scala 116:45]
      invalid_due_to_not_ready_i <= 1'h0; // @[cu_handler.scala 116:45]
    end else if (2'h1 == alloc_st) begin // @[cu_handler.scala 127:21]
      invalid_due_to_not_ready_i <= 1'h0; // @[cu_handler.scala 124:32]
    end else begin
      invalid_due_to_not_ready_i <= 2'h2 == alloc_st & _GEN_29;
    end
    if (reset) begin // @[cu_handler.scala 121:39]
      next_free_slot_valid <= 1'h0; // @[cu_handler.scala 121:39]
    end else begin
      next_free_slot_valid <= found_free_slot_valid2; // @[cu_handler.scala 122:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  next_free_slot = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  used_slot_bitmap_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  used_slot_bitmap_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  used_slot_bitmap_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  used_slot_bitmap_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pending_wg_bitmap_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pending_wg_bitmap_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pending_wg_bitmap_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pending_wg_bitmap_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pending_wf_count_0 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  pending_wf_count_1 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  pending_wf_count_2 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  pending_wf_count_3 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  curr_alloc_wf_count = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  curr_alloc_wf_slot = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  dispatch2cu_wf_dispatch_i = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dispatch2cu_wf_tag_dispatch_i = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  next_served_dealloc_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  next_served_dealloc = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  curr_dealloc_wg_slot = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  info_ram_rd_en = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  info_ram_rd_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  info_ram_wr_en = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  info_ram_wr_addr = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  info_ram_wr_reg = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  wg_done_valid_i = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  wg_done_wg_id_i = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  curr_wf_count = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  alloc_st = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  dealloc_st = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  invalid_due_to_not_ready_i = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  next_free_slot_valid = _RAND_31[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module gpu_interface(
  input         clock,
  input         reset,
  input         io_inflight_wg_buffer_gpu_valid,
  input  [9:0]  io_inflight_wg_buffer_gpu_wf_size,
  input  [31:0] io_inflight_wg_buffer_start_pc,
  input  [11:0] io_inflight_wg_buffer_gpu_vgpr_size_per_wf,
  input  [11:0] io_inflight_wg_buffer_gpu_sgpr_size_per_wf,
  input  [4:0]  io_allocator_wg_id_out,
  input  [1:0]  io_allocator_cu_id_out,
  input  [2:0]  io_allocator_wf_count,
  input  [11:0] io_allocator_vgpr_start_out,
  input  [11:0] io_allocator_sgpr_start_out,
  input  [11:0] io_allocator_lds_start_out,
  input         io_dis_controller_wg_alloc_valid,
  input         io_dis_controller_wg_dealloc_valid,
  output        io_gpu_interface_alloc_available,
  output        io_gpu_interface_dealloc_available,
  output [1:0]  io_gpu_interface_cu_id,
  output [4:0]  io_gpu_interface_dealloc_wg_id,
  output [1:0]  io_dispatch2cu_wf_dispatch,
  output [2:0]  io_dispatch2cu_wg_wf_count,
  output [9:0]  io_dispatch2cu_wf_size_dispatch,
  output [12:0] io_dispatch2cu_sgpr_base_dispatch,
  output [12:0] io_dispatch2cu_vgpr_base_dispatch,
  output [4:0]  io_dispatch2cu_wf_tag_dispatch,
  output [12:0] io_dispatch2cu_lds_base_dispatch,
  output [31:0] io_dispatch2cu_start_pc_dispatch,
  input  [1:0]  io_cu2dispatch_wf_done,
  input  [4:0]  io_cu2dispatch_wf_tag_done_0,
  input  [4:0]  io_cu2dispatch_wf_tag_done_1,
  input         io_cu2dispatch_ready_for_dispatch_0,
  input         io_cu2dispatch_ready_for_dispatch_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  wire  cu_handler_clock; // @[gpu_interface.scala 112:32]
  wire  cu_handler_reset; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_wg_alloc_en; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_io_wg_alloc_wg_id; // @[gpu_interface.scala 112:32]
  wire [2:0] cu_handler_io_wg_alloc_wf_count; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_ready_for_dispatch2cu; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_dispatch2cu_wf_dispatch; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_io_dispatch2cu_wf_tag_dispatch; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_cu2dispatch_wf_done_i; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_io_cu2dispatch_wf_tag_done_i; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_wg_done_ack; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_wg_done_valid; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_io_wg_done_wg_id; // @[gpu_interface.scala 112:32]
  wire  cu_handler_io_invalid_due_to_not_ready; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_clock; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_reset; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_wg_alloc_en; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_1_io_wg_alloc_wg_id; // @[gpu_interface.scala 112:32]
  wire [2:0] cu_handler_1_io_wg_alloc_wf_count; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_ready_for_dispatch2cu; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_dispatch2cu_wf_dispatch; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_1_io_dispatch2cu_wf_tag_dispatch; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_cu2dispatch_wf_done_i; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_1_io_cu2dispatch_wf_tag_done_i; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_wg_done_ack; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_wg_done_valid; // @[gpu_interface.scala 112:32]
  wire [4:0] cu_handler_1_io_wg_done_wg_id; // @[gpu_interface.scala 112:32]
  wire  cu_handler_1_io_invalid_due_to_not_ready; // @[gpu_interface.scala 112:32]
  reg  gpu_interface_dealloc_available_i; // @[gpu_interface.scala 46:52]
  reg  dis_controller_wg_dealloc_valid_i; // @[gpu_interface.scala 47:52]
  reg  handler_wg_done_ack_0; // @[gpu_interface.scala 48:38]
  reg  handler_wg_done_ack_1; // @[gpu_interface.scala 48:38]
  reg  chosen_done_cu_valid; // @[gpu_interface.scala 49:39]
  reg [1:0] chosen_done_cu_id; // @[gpu_interface.scala 51:36]
  reg  handler_wg_done_valid_0; // @[gpu_interface.scala 53:40]
  reg  handler_wg_done_valid_1; // @[gpu_interface.scala 53:40]
  reg [4:0] handler_wg_done_wg_id_0; // @[gpu_interface.scala 54:40]
  reg [4:0] handler_wg_done_wg_id_1; // @[gpu_interface.scala 54:40]
  reg  cu2dispatch_wf_done_i_0; // @[gpu_interface.scala 55:40]
  reg  cu2dispatch_wf_done_i_1; // @[gpu_interface.scala 55:40]
  reg [4:0] cu2dispatch_wf_tag_done_i_0; // @[gpu_interface.scala 56:44]
  reg [4:0] cu2dispatch_wf_tag_done_i_1; // @[gpu_interface.scala 56:44]
  reg [4:0] dealloc_st; // @[gpu_interface.scala 62:29]
  reg  dis_controller_wg_alloc_valid_i; // @[gpu_interface.scala 68:50]
  reg  inflight_wg_buffer_gpu_valid_i; // @[gpu_interface.scala 69:49]
  reg [9:0] inflight_wg_buffer_gpu_wf_size_i; // @[gpu_interface.scala 70:51]
  reg [31:0] inflight_wg_buffer_start_pc_i; // @[gpu_interface.scala 71:48]
  reg [11:0] inflight_wg_buffer_gpu_vgpr_size_per_wf_i; // @[gpu_interface.scala 72:60]
  reg [11:0] inflight_wg_buffer_gpu_sgpr_size_per_wf_i; // @[gpu_interface.scala 73:60]
  reg [4:0] allocator_wg_id_out_i; // @[gpu_interface.scala 75:40]
  reg [1:0] allocator_cu_id_out_i; // @[gpu_interface.scala 76:40]
  reg [2:0] allocator_wf_count_i; // @[gpu_interface.scala 77:39]
  reg [11:0] allocator_vgpr_start_out_i; // @[gpu_interface.scala 78:45]
  reg [11:0] allocator_sgpr_start_out_i; // @[gpu_interface.scala 79:45]
  reg [11:0] allocator_lds_start_out_i; // @[gpu_interface.scala 80:44]
  reg  gpu_interface_alloc_available_i; // @[gpu_interface.scala 82:50]
  reg [1:0] gpu_interface_cu_id_i; // @[gpu_interface.scala 83:40]
  reg [4:0] gpu_interface_dealloc_wg_id_i; // @[gpu_interface.scala 84:48]
  reg  dispatch2cu_wf_dispatch_handlers_0; // @[gpu_interface.scala 86:51]
  reg  dispatch2cu_wf_dispatch_handlers_1; // @[gpu_interface.scala 86:51]
  reg  invalid_due_to_not_ready_handlers_0; // @[gpu_interface.scala 87:52]
  reg  invalid_due_to_not_ready_handlers_1; // @[gpu_interface.scala 87:52]
  reg [4:0] dispatch2cu_wf_tag_dispatch_handlers_0; // @[gpu_interface.scala 88:55]
  reg [4:0] dispatch2cu_wf_tag_dispatch_handlers_1; // @[gpu_interface.scala 88:55]
  reg  handler_wg_alloc_en_0; // @[gpu_interface.scala 90:38]
  reg  handler_wg_alloc_en_1; // @[gpu_interface.scala 90:38]
  reg [4:0] handler_wg_alloc_wg_id_0; // @[gpu_interface.scala 91:41]
  reg [4:0] handler_wg_alloc_wg_id_1; // @[gpu_interface.scala 91:41]
  reg [2:0] handler_wg_alloc_wf_count_0; // @[gpu_interface.scala 92:44]
  reg [2:0] handler_wg_alloc_wf_count_1; // @[gpu_interface.scala 92:44]
  reg [1:0] dispatch2cu_wf_dispatch_i; // @[gpu_interface.scala 94:44]
  reg [2:0] dispatch2cu_wg_wf_count_i; // @[gpu_interface.scala 95:44]
  reg [9:0] dispatch2cu_wf_size_dispatch_i; // @[gpu_interface.scala 96:49]
  reg [12:0] dispatch2cu_sgpr_base_dispatch_i; // @[gpu_interface.scala 97:51]
  reg [12:0] dispatch2cu_vgpr_base_dispatch_i; // @[gpu_interface.scala 98:51]
  reg [4:0] dispatch2cu_wf_tag_dispatch_i; // @[gpu_interface.scala 99:48]
  reg [12:0] dispatch2cu_lds_base_dispatch_i; // @[gpu_interface.scala 100:50]
  reg [31:0] dispatch2cu_start_pc_dispatch_i; // @[gpu_interface.scala 101:50]
  reg [3:0] alloc_st; // @[gpu_interface.scala 108:27]
  wire  _GEN_10 = ~allocator_cu_id_out_i[0]; // @[gpu_interface.scala 146:25 154:{64,64}]
  wire [4:0] _GEN_12 = ~allocator_cu_id_out_i[0] ? allocator_wg_id_out_i : handler_wg_alloc_wg_id_0; // @[gpu_interface.scala 155:{67,67} 91:41]
  wire [4:0] _GEN_13 = allocator_cu_id_out_i[0] ? allocator_wg_id_out_i : handler_wg_alloc_wg_id_1; // @[gpu_interface.scala 155:{67,67} 91:41]
  wire [2:0] _GEN_14 = ~allocator_cu_id_out_i[0] ? allocator_wf_count_i : handler_wg_alloc_wf_count_0; // @[gpu_interface.scala 156:{70,70} 92:44]
  wire [2:0] _GEN_15 = allocator_cu_id_out_i[0] ? allocator_wf_count_i : handler_wg_alloc_wf_count_1; // @[gpu_interface.scala 156:{70,70} 92:44]
  wire  _GEN_16 = inflight_wg_buffer_gpu_valid_i & _GEN_10; // @[gpu_interface.scala 146:25 153:53]
  wire  _GEN_17 = inflight_wg_buffer_gpu_valid_i & allocator_cu_id_out_i[0]; // @[gpu_interface.scala 146:25 153:53]
  wire [4:0] _GEN_18 = inflight_wg_buffer_gpu_valid_i ? _GEN_12 : handler_wg_alloc_wg_id_0; // @[gpu_interface.scala 153:53 91:41]
  wire [4:0] _GEN_19 = inflight_wg_buffer_gpu_valid_i ? _GEN_13 : handler_wg_alloc_wg_id_1; // @[gpu_interface.scala 153:53 91:41]
  wire [2:0] _GEN_20 = inflight_wg_buffer_gpu_valid_i ? _GEN_14 : handler_wg_alloc_wf_count_0; // @[gpu_interface.scala 153:53 92:44]
  wire [2:0] _GEN_21 = inflight_wg_buffer_gpu_valid_i ? _GEN_15 : handler_wg_alloc_wf_count_1; // @[gpu_interface.scala 153:53 92:44]
  wire [2:0] _GEN_23 = inflight_wg_buffer_gpu_valid_i ? 3'h4 : 3'h2; // @[gpu_interface.scala 153:53 158:30 162:30]
  wire  _GEN_24 = dis_controller_wg_alloc_valid_i & _GEN_16; // @[gpu_interface.scala 146:25 152:50]
  wire  _GEN_25 = dis_controller_wg_alloc_valid_i & _GEN_17; // @[gpu_interface.scala 146:25 152:50]
  wire  _GEN_47 = allocator_cu_id_out_i[0] ? dispatch2cu_wf_dispatch_handlers_1 : dispatch2cu_wf_dispatch_handlers_0; // @[gpu_interface.scala 176:{74,74}]
  wire [3:0] _dispatch2cu_wf_dispatch_i_T = 4'h1 << allocator_cu_id_out_i; // @[gpu_interface.scala 177:50]
  wire [4:0] _GEN_49 = allocator_cu_id_out_i[0] ? dispatch2cu_wf_tag_dispatch_handlers_1 :
    dispatch2cu_wf_tag_dispatch_handlers_0; // @[gpu_interface.scala 178:{47,47}]
  wire [3:0] _GEN_50 = _GEN_47 ? _dispatch2cu_wf_dispatch_i_T : 4'h0; // @[gpu_interface.scala 147:31 176:74 177:43]
  wire [4:0] _GEN_51 = _GEN_47 ? _GEN_49 : dispatch2cu_wf_tag_dispatch_i; // @[gpu_interface.scala 176:74 178:47 99:48]
  wire [2:0] _GEN_52 = _GEN_47 ? allocator_wf_count_i : dispatch2cu_wg_wf_count_i; // @[gpu_interface.scala 176:74 179:43 95:44]
  wire [9:0] _GEN_53 = _GEN_47 ? inflight_wg_buffer_gpu_wf_size_i : dispatch2cu_wf_size_dispatch_i; // @[gpu_interface.scala 176:74 181:48 96:49]
  wire [31:0] _GEN_54 = _GEN_47 ? inflight_wg_buffer_start_pc_i : dispatch2cu_start_pc_dispatch_i; // @[gpu_interface.scala 176:74 182:49 101:50]
  wire [12:0] _GEN_55 = _GEN_47 ? {{1'd0}, allocator_vgpr_start_out_i} : dispatch2cu_vgpr_base_dispatch_i; // @[gpu_interface.scala 176:74 183:50 98:51]
  wire [12:0] _GEN_56 = _GEN_47 ? {{1'd0}, allocator_sgpr_start_out_i} : dispatch2cu_sgpr_base_dispatch_i; // @[gpu_interface.scala 176:74 184:50 97:51]
  wire [12:0] _GEN_57 = _GEN_47 ? {{1'd0}, allocator_lds_start_out_i} : dispatch2cu_lds_base_dispatch_i; // @[gpu_interface.scala 176:74 185:49 100:50]
  wire [3:0] _GEN_58 = _GEN_47 ? 4'h8 : alloc_st; // @[gpu_interface.scala 176:74 186:26 108:27]
  wire [12:0] _GEN_145 = {{1'd0}, inflight_wg_buffer_gpu_sgpr_size_per_wf_i}; // @[gpu_interface.scala 193:86]
  wire [12:0] _dispatch2cu_sgpr_base_dispatch_i_T_1 = dispatch2cu_sgpr_base_dispatch_i + _GEN_145; // @[gpu_interface.scala 193:86]
  wire [12:0] _GEN_146 = {{1'd0}, inflight_wg_buffer_gpu_vgpr_size_per_wf_i}; // @[gpu_interface.scala 194:86]
  wire [12:0] _dispatch2cu_vgpr_base_dispatch_i_T_1 = dispatch2cu_vgpr_base_dispatch_i + _GEN_146; // @[gpu_interface.scala 194:86]
  wire  _GEN_64 = allocator_cu_id_out_i[0] ? invalid_due_to_not_ready_handlers_1 : invalid_due_to_not_ready_handlers_0; // @[gpu_interface.scala 196:{80,80}]
  wire  _GEN_66 = _GEN_64 ? gpu_interface_alloc_available_i : 1'h1; // @[gpu_interface.scala 196:80 200:49 82:50]
  wire [3:0] _GEN_67 = _GEN_64 ? alloc_st : 4'h1; // @[gpu_interface.scala 108:27 196:80 201:26]
  wire [12:0] _GEN_70 = _GEN_47 ? _dispatch2cu_sgpr_base_dispatch_i_T_1 : dispatch2cu_sgpr_base_dispatch_i; // @[gpu_interface.scala 190:74 193:50 97:51]
  wire [12:0] _GEN_71 = _GEN_47 ? _dispatch2cu_vgpr_base_dispatch_i_T_1 : dispatch2cu_vgpr_base_dispatch_i; // @[gpu_interface.scala 190:74 194:50 98:51]
  wire  _GEN_72 = _GEN_47 ? gpu_interface_alloc_available_i : _GEN_66; // @[gpu_interface.scala 190:74 82:50]
  wire [3:0] _GEN_73 = _GEN_47 ? alloc_st : _GEN_67; // @[gpu_interface.scala 108:27 190:74]
  wire [3:0] _GEN_74 = 4'h8 == alloc_st ? _GEN_50 : 4'h0; // @[gpu_interface.scala 149:21 147:31]
  wire [4:0] _GEN_75 = 4'h8 == alloc_st ? _GEN_51 : dispatch2cu_wf_tag_dispatch_i; // @[gpu_interface.scala 149:21 99:48]
  wire [12:0] _GEN_76 = 4'h8 == alloc_st ? _GEN_70 : dispatch2cu_sgpr_base_dispatch_i; // @[gpu_interface.scala 149:21 97:51]
  wire [12:0] _GEN_77 = 4'h8 == alloc_st ? _GEN_71 : dispatch2cu_vgpr_base_dispatch_i; // @[gpu_interface.scala 149:21 98:51]
  wire  _GEN_78 = 4'h8 == alloc_st ? _GEN_72 : gpu_interface_alloc_available_i; // @[gpu_interface.scala 149:21 82:50]
  wire [3:0] _GEN_79 = 4'h8 == alloc_st ? _GEN_73 : alloc_st; // @[gpu_interface.scala 149:21 108:27]
  wire [3:0] _GEN_80 = 4'h4 == alloc_st ? _GEN_50 : _GEN_74; // @[gpu_interface.scala 149:21]
  wire  _GEN_90 = 4'h2 == alloc_st & _GEN_16; // @[gpu_interface.scala 149:21 146:25]
  wire  _GEN_91 = 4'h2 == alloc_st & _GEN_17; // @[gpu_interface.scala 149:21 146:25]
  wire [3:0] _GEN_98 = 4'h2 == alloc_st ? 4'h0 : _GEN_80; // @[gpu_interface.scala 149:21 147:31]
  wire [3:0] _GEN_114 = 4'h1 == alloc_st ? 4'h0 : _GEN_98; // @[gpu_interface.scala 149:21 147:31]
  wire  _GEN_122 = ~chosen_done_cu_id[0]; // @[gpu_interface.scala 219:25 227:{56,56}]
  wire  _GEN_128 = chosen_done_cu_valid & _GEN_122; // @[gpu_interface.scala 219:25 224:39]
  wire  _GEN_129 = chosen_done_cu_valid & chosen_done_cu_id[0]; // @[gpu_interface.scala 219:25 224:39]
  wire  _GEN_133 = dis_controller_wg_dealloc_valid_i ? 1'h0 : 1'h1; // @[gpu_interface.scala 218:39 233:52 237:51]
  wire  _GEN_135 = 5'h2 == dealloc_st & _GEN_133; // @[gpu_interface.scala 222:23 218:39]
  wire  _GEN_138 = 5'h1 == dealloc_st & _GEN_128; // @[gpu_interface.scala 222:23 219:25]
  wire  _GEN_139 = 5'h1 == dealloc_st & _GEN_129; // @[gpu_interface.scala 222:23 219:25]
  wire  cu_found_valid = handler_wg_done_valid_0 | handler_wg_done_valid_1; // @[gpu_interface.scala 247:39 248:28]
  wire  _GEN_144 = handler_wg_done_valid_0 ? 1'h0 : handler_wg_done_valid_1; // @[gpu_interface.scala 247:39 249:22]
  wire [1:0] cu_found = {{1'd0}, _GEN_144}; // @[gpu_interface.scala 243:24]
  wire [3:0] _GEN_147 = reset ? 4'h0 : _GEN_114; // @[gpu_interface.scala 94:{44,44}]
  cu_handler cu_handler ( // @[gpu_interface.scala 112:32]
    .clock(cu_handler_clock),
    .reset(cu_handler_reset),
    .io_wg_alloc_en(cu_handler_io_wg_alloc_en),
    .io_wg_alloc_wg_id(cu_handler_io_wg_alloc_wg_id),
    .io_wg_alloc_wf_count(cu_handler_io_wg_alloc_wf_count),
    .io_ready_for_dispatch2cu(cu_handler_io_ready_for_dispatch2cu),
    .io_dispatch2cu_wf_dispatch(cu_handler_io_dispatch2cu_wf_dispatch),
    .io_dispatch2cu_wf_tag_dispatch(cu_handler_io_dispatch2cu_wf_tag_dispatch),
    .io_cu2dispatch_wf_done_i(cu_handler_io_cu2dispatch_wf_done_i),
    .io_cu2dispatch_wf_tag_done_i(cu_handler_io_cu2dispatch_wf_tag_done_i),
    .io_wg_done_ack(cu_handler_io_wg_done_ack),
    .io_wg_done_valid(cu_handler_io_wg_done_valid),
    .io_wg_done_wg_id(cu_handler_io_wg_done_wg_id),
    .io_invalid_due_to_not_ready(cu_handler_io_invalid_due_to_not_ready)
  );
  cu_handler cu_handler_1 ( // @[gpu_interface.scala 112:32]
    .clock(cu_handler_1_clock),
    .reset(cu_handler_1_reset),
    .io_wg_alloc_en(cu_handler_1_io_wg_alloc_en),
    .io_wg_alloc_wg_id(cu_handler_1_io_wg_alloc_wg_id),
    .io_wg_alloc_wf_count(cu_handler_1_io_wg_alloc_wf_count),
    .io_ready_for_dispatch2cu(cu_handler_1_io_ready_for_dispatch2cu),
    .io_dispatch2cu_wf_dispatch(cu_handler_1_io_dispatch2cu_wf_dispatch),
    .io_dispatch2cu_wf_tag_dispatch(cu_handler_1_io_dispatch2cu_wf_tag_dispatch),
    .io_cu2dispatch_wf_done_i(cu_handler_1_io_cu2dispatch_wf_done_i),
    .io_cu2dispatch_wf_tag_done_i(cu_handler_1_io_cu2dispatch_wf_tag_done_i),
    .io_wg_done_ack(cu_handler_1_io_wg_done_ack),
    .io_wg_done_valid(cu_handler_1_io_wg_done_valid),
    .io_wg_done_wg_id(cu_handler_1_io_wg_done_wg_id),
    .io_invalid_due_to_not_ready(cu_handler_1_io_invalid_due_to_not_ready)
  );
  assign io_gpu_interface_alloc_available = gpu_interface_alloc_available_i; // @[gpu_interface.scala 257:38]
  assign io_gpu_interface_dealloc_available = gpu_interface_dealloc_available_i; // @[gpu_interface.scala 254:40]
  assign io_gpu_interface_cu_id = gpu_interface_cu_id_i; // @[gpu_interface.scala 256:28]
  assign io_gpu_interface_dealloc_wg_id = gpu_interface_dealloc_wg_id_i; // @[gpu_interface.scala 255:36]
  assign io_dispatch2cu_wf_dispatch = dispatch2cu_wf_dispatch_i; // @[gpu_interface.scala 258:32]
  assign io_dispatch2cu_wg_wf_count = dispatch2cu_wg_wf_count_i; // @[gpu_interface.scala 260:32]
  assign io_dispatch2cu_wf_size_dispatch = dispatch2cu_wf_size_dispatch_i; // @[gpu_interface.scala 261:37]
  assign io_dispatch2cu_sgpr_base_dispatch = dispatch2cu_sgpr_base_dispatch_i; // @[gpu_interface.scala 262:39]
  assign io_dispatch2cu_vgpr_base_dispatch = dispatch2cu_vgpr_base_dispatch_i; // @[gpu_interface.scala 263:39]
  assign io_dispatch2cu_wf_tag_dispatch = dispatch2cu_wf_tag_dispatch_i; // @[gpu_interface.scala 259:36]
  assign io_dispatch2cu_lds_base_dispatch = dispatch2cu_lds_base_dispatch_i; // @[gpu_interface.scala 264:38]
  assign io_dispatch2cu_start_pc_dispatch = dispatch2cu_start_pc_dispatch_i; // @[gpu_interface.scala 265:38]
  assign cu_handler_clock = clock;
  assign cu_handler_reset = reset;
  assign cu_handler_io_wg_alloc_en = handler_wg_alloc_en_0; // @[gpu_interface.scala 113:35]
  assign cu_handler_io_wg_alloc_wg_id = handler_wg_alloc_wg_id_0; // @[gpu_interface.scala 114:38]
  assign cu_handler_io_wg_alloc_wf_count = handler_wg_alloc_wf_count_0; // @[gpu_interface.scala 115:41]
  assign cu_handler_io_ready_for_dispatch2cu = io_cu2dispatch_ready_for_dispatch_0; // @[gpu_interface.scala 119:45]
  assign cu_handler_io_cu2dispatch_wf_done_i = cu2dispatch_wf_done_i_0; // @[gpu_interface.scala 116:45]
  assign cu_handler_io_cu2dispatch_wf_tag_done_i = cu2dispatch_wf_tag_done_i_0; // @[gpu_interface.scala 117:49]
  assign cu_handler_io_wg_done_ack = handler_wg_done_ack_0; // @[gpu_interface.scala 118:35]
  assign cu_handler_1_clock = clock;
  assign cu_handler_1_reset = reset;
  assign cu_handler_1_io_wg_alloc_en = handler_wg_alloc_en_1; // @[gpu_interface.scala 113:35]
  assign cu_handler_1_io_wg_alloc_wg_id = handler_wg_alloc_wg_id_1; // @[gpu_interface.scala 114:38]
  assign cu_handler_1_io_wg_alloc_wf_count = handler_wg_alloc_wf_count_1; // @[gpu_interface.scala 115:41]
  assign cu_handler_1_io_ready_for_dispatch2cu = io_cu2dispatch_ready_for_dispatch_1; // @[gpu_interface.scala 119:45]
  assign cu_handler_1_io_cu2dispatch_wf_done_i = cu2dispatch_wf_done_i_1; // @[gpu_interface.scala 116:45]
  assign cu_handler_1_io_cu2dispatch_wf_tag_done_i = cu2dispatch_wf_tag_done_i_1; // @[gpu_interface.scala 117:49]
  assign cu_handler_1_io_wg_done_ack = handler_wg_done_ack_1; // @[gpu_interface.scala 118:35]
  always @(posedge clock) begin
    if (reset) begin // @[gpu_interface.scala 46:52]
      gpu_interface_dealloc_available_i <= 1'h0; // @[gpu_interface.scala 46:52]
    end else if (5'h1 == dealloc_st) begin // @[gpu_interface.scala 222:23]
      gpu_interface_dealloc_available_i <= chosen_done_cu_valid;
    end else begin
      gpu_interface_dealloc_available_i <= _GEN_135;
    end
    if (reset) begin // @[gpu_interface.scala 47:52]
      dis_controller_wg_dealloc_valid_i <= 1'h0; // @[gpu_interface.scala 47:52]
    end else begin
      dis_controller_wg_dealloc_valid_i <= io_dis_controller_wg_dealloc_valid; // @[gpu_interface.scala 214:39]
    end
    if (reset) begin // @[gpu_interface.scala 48:38]
      handler_wg_done_ack_0 <= 1'h0; // @[gpu_interface.scala 48:38]
    end else begin
      handler_wg_done_ack_0 <= _GEN_138;
    end
    if (reset) begin // @[gpu_interface.scala 48:38]
      handler_wg_done_ack_1 <= 1'h0; // @[gpu_interface.scala 48:38]
    end else begin
      handler_wg_done_ack_1 <= _GEN_139;
    end
    if (reset) begin // @[gpu_interface.scala 49:39]
      chosen_done_cu_valid <= 1'h0; // @[gpu_interface.scala 49:39]
    end else begin
      chosen_done_cu_valid <= cu_found_valid; // @[gpu_interface.scala 215:26]
    end
    if (reset) begin // @[gpu_interface.scala 51:36]
      chosen_done_cu_id <= 2'h0; // @[gpu_interface.scala 51:36]
    end else begin
      chosen_done_cu_id <= cu_found; // @[gpu_interface.scala 216:23]
    end
    if (reset) begin // @[gpu_interface.scala 53:40]
      handler_wg_done_valid_0 <= 1'h0; // @[gpu_interface.scala 53:40]
    end else begin
      handler_wg_done_valid_0 <= cu_handler_io_wg_done_valid; // @[gpu_interface.scala 122:34]
    end
    if (reset) begin // @[gpu_interface.scala 53:40]
      handler_wg_done_valid_1 <= 1'h0; // @[gpu_interface.scala 53:40]
    end else begin
      handler_wg_done_valid_1 <= cu_handler_1_io_wg_done_valid; // @[gpu_interface.scala 122:34]
    end
    if (reset) begin // @[gpu_interface.scala 54:40]
      handler_wg_done_wg_id_0 <= 5'h0; // @[gpu_interface.scala 54:40]
    end else begin
      handler_wg_done_wg_id_0 <= cu_handler_io_wg_done_wg_id; // @[gpu_interface.scala 123:34]
    end
    if (reset) begin // @[gpu_interface.scala 54:40]
      handler_wg_done_wg_id_1 <= 5'h0; // @[gpu_interface.scala 54:40]
    end else begin
      handler_wg_done_wg_id_1 <= cu_handler_1_io_wg_done_wg_id; // @[gpu_interface.scala 123:34]
    end
    if (reset) begin // @[gpu_interface.scala 55:40]
      cu2dispatch_wf_done_i_0 <= 1'h0; // @[gpu_interface.scala 55:40]
    end else begin
      cu2dispatch_wf_done_i_0 <= io_cu2dispatch_wf_done[0]; // @[gpu_interface.scala 205:27]
    end
    if (reset) begin // @[gpu_interface.scala 55:40]
      cu2dispatch_wf_done_i_1 <= 1'h0; // @[gpu_interface.scala 55:40]
    end else begin
      cu2dispatch_wf_done_i_1 <= io_cu2dispatch_wf_done[1]; // @[gpu_interface.scala 205:27]
    end
    if (reset) begin // @[gpu_interface.scala 56:44]
      cu2dispatch_wf_tag_done_i_0 <= 5'h0; // @[gpu_interface.scala 56:44]
    end else begin
      cu2dispatch_wf_tag_done_i_0 <= io_cu2dispatch_wf_tag_done_0; // @[gpu_interface.scala 208:38]
    end
    if (reset) begin // @[gpu_interface.scala 56:44]
      cu2dispatch_wf_tag_done_i_1 <= 5'h0; // @[gpu_interface.scala 56:44]
    end else begin
      cu2dispatch_wf_tag_done_i_1 <= io_cu2dispatch_wf_tag_done_1; // @[gpu_interface.scala 208:38]
    end
    if (reset) begin // @[gpu_interface.scala 62:29]
      dealloc_st <= 5'h1; // @[gpu_interface.scala 62:29]
    end else if (5'h1 == dealloc_st) begin // @[gpu_interface.scala 222:23]
      if (chosen_done_cu_valid) begin // @[gpu_interface.scala 224:39]
        dealloc_st <= 5'h2; // @[gpu_interface.scala 229:28]
      end
    end else if (5'h2 == dealloc_st) begin // @[gpu_interface.scala 222:23]
      if (dis_controller_wg_dealloc_valid_i) begin // @[gpu_interface.scala 233:52]
        dealloc_st <= 5'h1; // @[gpu_interface.scala 234:28]
      end
    end
    if (reset) begin // @[gpu_interface.scala 68:50]
      dis_controller_wg_alloc_valid_i <= 1'h0; // @[gpu_interface.scala 68:50]
    end else begin
      dis_controller_wg_alloc_valid_i <= io_dis_controller_wg_alloc_valid; // @[gpu_interface.scala 126:37]
    end
    if (reset) begin // @[gpu_interface.scala 69:49]
      inflight_wg_buffer_gpu_valid_i <= 1'h0; // @[gpu_interface.scala 69:49]
    end else begin
      inflight_wg_buffer_gpu_valid_i <= io_inflight_wg_buffer_gpu_valid; // @[gpu_interface.scala 127:36]
    end
    if (reset) begin // @[gpu_interface.scala 70:51]
      inflight_wg_buffer_gpu_wf_size_i <= 10'h0; // @[gpu_interface.scala 70:51]
    end else if (io_inflight_wg_buffer_gpu_valid) begin // @[gpu_interface.scala 128:42]
      inflight_wg_buffer_gpu_wf_size_i <= io_inflight_wg_buffer_gpu_wf_size; // @[gpu_interface.scala 129:42]
    end
    if (reset) begin // @[gpu_interface.scala 71:48]
      inflight_wg_buffer_start_pc_i <= 32'h0; // @[gpu_interface.scala 71:48]
    end else if (io_inflight_wg_buffer_gpu_valid) begin // @[gpu_interface.scala 128:42]
      inflight_wg_buffer_start_pc_i <= io_inflight_wg_buffer_start_pc; // @[gpu_interface.scala 130:39]
    end
    if (reset) begin // @[gpu_interface.scala 72:60]
      inflight_wg_buffer_gpu_vgpr_size_per_wf_i <= 12'h0; // @[gpu_interface.scala 72:60]
    end else if (io_inflight_wg_buffer_gpu_valid) begin // @[gpu_interface.scala 128:42]
      inflight_wg_buffer_gpu_vgpr_size_per_wf_i <= io_inflight_wg_buffer_gpu_vgpr_size_per_wf; // @[gpu_interface.scala 131:51]
    end
    if (reset) begin // @[gpu_interface.scala 73:60]
      inflight_wg_buffer_gpu_sgpr_size_per_wf_i <= 12'h0; // @[gpu_interface.scala 73:60]
    end else if (io_inflight_wg_buffer_gpu_valid) begin // @[gpu_interface.scala 128:42]
      inflight_wg_buffer_gpu_sgpr_size_per_wf_i <= io_inflight_wg_buffer_gpu_sgpr_size_per_wf; // @[gpu_interface.scala 132:51]
    end
    if (reset) begin // @[gpu_interface.scala 75:40]
      allocator_wg_id_out_i <= 5'h0; // @[gpu_interface.scala 75:40]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[gpu_interface.scala 134:43]
      allocator_wg_id_out_i <= io_allocator_wg_id_out; // @[gpu_interface.scala 135:31]
    end
    if (reset) begin // @[gpu_interface.scala 76:40]
      allocator_cu_id_out_i <= 2'h0; // @[gpu_interface.scala 76:40]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[gpu_interface.scala 134:43]
      allocator_cu_id_out_i <= io_allocator_cu_id_out; // @[gpu_interface.scala 136:31]
    end
    if (reset) begin // @[gpu_interface.scala 77:39]
      allocator_wf_count_i <= 3'h0; // @[gpu_interface.scala 77:39]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[gpu_interface.scala 134:43]
      allocator_wf_count_i <= io_allocator_wf_count; // @[gpu_interface.scala 137:30]
    end
    if (reset) begin // @[gpu_interface.scala 78:45]
      allocator_vgpr_start_out_i <= 12'h0; // @[gpu_interface.scala 78:45]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[gpu_interface.scala 134:43]
      allocator_vgpr_start_out_i <= io_allocator_vgpr_start_out; // @[gpu_interface.scala 138:36]
    end
    if (reset) begin // @[gpu_interface.scala 79:45]
      allocator_sgpr_start_out_i <= 12'h0; // @[gpu_interface.scala 79:45]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[gpu_interface.scala 134:43]
      allocator_sgpr_start_out_i <= io_allocator_sgpr_start_out; // @[gpu_interface.scala 139:36]
    end
    if (reset) begin // @[gpu_interface.scala 80:44]
      allocator_lds_start_out_i <= 12'h0; // @[gpu_interface.scala 80:44]
    end else if (io_dis_controller_wg_alloc_valid) begin // @[gpu_interface.scala 134:43]
      allocator_lds_start_out_i <= io_allocator_lds_start_out; // @[gpu_interface.scala 140:35]
    end
    if (reset) begin // @[gpu_interface.scala 82:50]
      gpu_interface_alloc_available_i <= 1'h0; // @[gpu_interface.scala 82:50]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (dis_controller_wg_alloc_valid_i) begin // @[gpu_interface.scala 152:50]
        gpu_interface_alloc_available_i <= 1'h0;
      end else begin
        gpu_interface_alloc_available_i <= 1'h1; // @[gpu_interface.scala 151:45]
      end
    end else if (4'h2 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (inflight_wg_buffer_gpu_valid_i) begin // @[gpu_interface.scala 167:49]
        gpu_interface_alloc_available_i <= 1'h0; // @[gpu_interface.scala 171:49]
      end
    end else if (!(4'h4 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      gpu_interface_alloc_available_i <= _GEN_78;
    end
    if (reset) begin // @[gpu_interface.scala 83:40]
      gpu_interface_cu_id_i <= 2'h0; // @[gpu_interface.scala 83:40]
    end else if (5'h1 == dealloc_st) begin // @[gpu_interface.scala 222:23]
      if (chosen_done_cu_valid) begin // @[gpu_interface.scala 224:39]
        gpu_interface_cu_id_i <= chosen_done_cu_id; // @[gpu_interface.scala 226:39]
      end
    end
    if (reset) begin // @[gpu_interface.scala 84:48]
      gpu_interface_dealloc_wg_id_i <= 5'h0; // @[gpu_interface.scala 84:48]
    end else if (5'h1 == dealloc_st) begin // @[gpu_interface.scala 222:23]
      if (chosen_done_cu_valid) begin // @[gpu_interface.scala 224:39]
        if (chosen_done_cu_id[0]) begin // @[gpu_interface.scala 228:47]
          gpu_interface_dealloc_wg_id_i <= handler_wg_done_wg_id_1; // @[gpu_interface.scala 228:47]
        end else begin
          gpu_interface_dealloc_wg_id_i <= handler_wg_done_wg_id_0;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 86:51]
      dispatch2cu_wf_dispatch_handlers_0 <= 1'h0; // @[gpu_interface.scala 86:51]
    end else begin
      dispatch2cu_wf_dispatch_handlers_0 <= cu_handler_io_dispatch2cu_wf_dispatch; // @[gpu_interface.scala 120:45]
    end
    if (reset) begin // @[gpu_interface.scala 86:51]
      dispatch2cu_wf_dispatch_handlers_1 <= 1'h0; // @[gpu_interface.scala 86:51]
    end else begin
      dispatch2cu_wf_dispatch_handlers_1 <= cu_handler_1_io_dispatch2cu_wf_dispatch; // @[gpu_interface.scala 120:45]
    end
    if (reset) begin // @[gpu_interface.scala 87:52]
      invalid_due_to_not_ready_handlers_0 <= 1'h0; // @[gpu_interface.scala 87:52]
    end else begin
      invalid_due_to_not_ready_handlers_0 <= cu_handler_io_invalid_due_to_not_ready; // @[gpu_interface.scala 124:46]
    end
    if (reset) begin // @[gpu_interface.scala 87:52]
      invalid_due_to_not_ready_handlers_1 <= 1'h0; // @[gpu_interface.scala 87:52]
    end else begin
      invalid_due_to_not_ready_handlers_1 <= cu_handler_1_io_invalid_due_to_not_ready; // @[gpu_interface.scala 124:46]
    end
    if (reset) begin // @[gpu_interface.scala 88:55]
      dispatch2cu_wf_tag_dispatch_handlers_0 <= 5'h0; // @[gpu_interface.scala 88:55]
    end else begin
      dispatch2cu_wf_tag_dispatch_handlers_0 <= cu_handler_io_dispatch2cu_wf_tag_dispatch; // @[gpu_interface.scala 121:49]
    end
    if (reset) begin // @[gpu_interface.scala 88:55]
      dispatch2cu_wf_tag_dispatch_handlers_1 <= 5'h0; // @[gpu_interface.scala 88:55]
    end else begin
      dispatch2cu_wf_tag_dispatch_handlers_1 <= cu_handler_1_io_dispatch2cu_wf_tag_dispatch; // @[gpu_interface.scala 121:49]
    end
    if (reset) begin // @[gpu_interface.scala 90:38]
      handler_wg_alloc_en_0 <= 1'h0; // @[gpu_interface.scala 90:38]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      handler_wg_alloc_en_0 <= _GEN_24;
    end else begin
      handler_wg_alloc_en_0 <= _GEN_90;
    end
    if (reset) begin // @[gpu_interface.scala 90:38]
      handler_wg_alloc_en_1 <= 1'h0; // @[gpu_interface.scala 90:38]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      handler_wg_alloc_en_1 <= _GEN_25;
    end else begin
      handler_wg_alloc_en_1 <= _GEN_91;
    end
    if (reset) begin // @[gpu_interface.scala 91:41]
      handler_wg_alloc_wg_id_0 <= 5'h0; // @[gpu_interface.scala 91:41]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (dis_controller_wg_alloc_valid_i) begin // @[gpu_interface.scala 152:50]
        handler_wg_alloc_wg_id_0 <= _GEN_18;
      end
    end else if (4'h2 == alloc_st) begin // @[gpu_interface.scala 149:21]
      handler_wg_alloc_wg_id_0 <= _GEN_18;
    end
    if (reset) begin // @[gpu_interface.scala 91:41]
      handler_wg_alloc_wg_id_1 <= 5'h0; // @[gpu_interface.scala 91:41]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (dis_controller_wg_alloc_valid_i) begin // @[gpu_interface.scala 152:50]
        handler_wg_alloc_wg_id_1 <= _GEN_19;
      end
    end else if (4'h2 == alloc_st) begin // @[gpu_interface.scala 149:21]
      handler_wg_alloc_wg_id_1 <= _GEN_19;
    end
    if (reset) begin // @[gpu_interface.scala 92:44]
      handler_wg_alloc_wf_count_0 <= 3'h0; // @[gpu_interface.scala 92:44]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (dis_controller_wg_alloc_valid_i) begin // @[gpu_interface.scala 152:50]
        handler_wg_alloc_wf_count_0 <= _GEN_20;
      end
    end else if (4'h2 == alloc_st) begin // @[gpu_interface.scala 149:21]
      handler_wg_alloc_wf_count_0 <= _GEN_20;
    end
    if (reset) begin // @[gpu_interface.scala 92:44]
      handler_wg_alloc_wf_count_1 <= 3'h0; // @[gpu_interface.scala 92:44]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (dis_controller_wg_alloc_valid_i) begin // @[gpu_interface.scala 152:50]
        handler_wg_alloc_wf_count_1 <= _GEN_21;
      end
    end else if (4'h2 == alloc_st) begin // @[gpu_interface.scala 149:21]
      handler_wg_alloc_wf_count_1 <= _GEN_21;
    end
    dispatch2cu_wf_dispatch_i <= _GEN_147[1:0]; // @[gpu_interface.scala 94:{44,44}]
    if (reset) begin // @[gpu_interface.scala 95:44]
      dispatch2cu_wg_wf_count_i <= 3'h0; // @[gpu_interface.scala 95:44]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_wg_wf_count_i <= _GEN_52;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 96:49]
      dispatch2cu_wf_size_dispatch_i <= 10'h0; // @[gpu_interface.scala 96:49]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_wf_size_dispatch_i <= _GEN_53;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 97:51]
      dispatch2cu_sgpr_base_dispatch_i <= 13'h0; // @[gpu_interface.scala 97:51]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_sgpr_base_dispatch_i <= _GEN_56;
        end else begin
          dispatch2cu_sgpr_base_dispatch_i <= _GEN_76;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 98:51]
      dispatch2cu_vgpr_base_dispatch_i <= 13'h0; // @[gpu_interface.scala 98:51]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_vgpr_base_dispatch_i <= _GEN_55;
        end else begin
          dispatch2cu_vgpr_base_dispatch_i <= _GEN_77;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 99:48]
      dispatch2cu_wf_tag_dispatch_i <= 5'h0; // @[gpu_interface.scala 99:48]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_wf_tag_dispatch_i <= _GEN_51;
        end else begin
          dispatch2cu_wf_tag_dispatch_i <= _GEN_75;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 100:50]
      dispatch2cu_lds_base_dispatch_i <= 13'h0; // @[gpu_interface.scala 100:50]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_lds_base_dispatch_i <= _GEN_57;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 101:50]
      dispatch2cu_start_pc_dispatch_i <= 32'h0; // @[gpu_interface.scala 101:50]
    end else if (!(4'h1 == alloc_st)) begin // @[gpu_interface.scala 149:21]
      if (!(4'h2 == alloc_st)) begin // @[gpu_interface.scala 149:21]
        if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
          dispatch2cu_start_pc_dispatch_i <= _GEN_54;
        end
      end
    end
    if (reset) begin // @[gpu_interface.scala 108:27]
      alloc_st <= 4'h1; // @[gpu_interface.scala 108:27]
    end else if (4'h1 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (dis_controller_wg_alloc_valid_i) begin // @[gpu_interface.scala 152:50]
        alloc_st <= {{1'd0}, _GEN_23};
      end
    end else if (4'h2 == alloc_st) begin // @[gpu_interface.scala 149:21]
      if (inflight_wg_buffer_gpu_valid_i) begin // @[gpu_interface.scala 167:49]
        alloc_st <= 4'h4; // @[gpu_interface.scala 172:26]
      end
    end else if (4'h4 == alloc_st) begin // @[gpu_interface.scala 149:21]
      alloc_st <= _GEN_58;
    end else begin
      alloc_st <= _GEN_79;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  gpu_interface_dealloc_available_i = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dis_controller_wg_dealloc_valid_i = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  handler_wg_done_ack_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  handler_wg_done_ack_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  chosen_done_cu_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  chosen_done_cu_id = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  handler_wg_done_valid_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  handler_wg_done_valid_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  handler_wg_done_wg_id_0 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  handler_wg_done_wg_id_1 = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  cu2dispatch_wf_done_i_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cu2dispatch_wf_done_i_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cu2dispatch_wf_tag_done_i_0 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  cu2dispatch_wf_tag_done_i_1 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  dealloc_st = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  dis_controller_wg_alloc_valid_i = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_valid_i = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_wf_size_i = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  inflight_wg_buffer_start_pc_i = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_vgpr_size_per_wf_i = _RAND_19[11:0];
  _RAND_20 = {1{`RANDOM}};
  inflight_wg_buffer_gpu_sgpr_size_per_wf_i = _RAND_20[11:0];
  _RAND_21 = {1{`RANDOM}};
  allocator_wg_id_out_i = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  allocator_cu_id_out_i = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  allocator_wf_count_i = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  allocator_vgpr_start_out_i = _RAND_24[11:0];
  _RAND_25 = {1{`RANDOM}};
  allocator_sgpr_start_out_i = _RAND_25[11:0];
  _RAND_26 = {1{`RANDOM}};
  allocator_lds_start_out_i = _RAND_26[11:0];
  _RAND_27 = {1{`RANDOM}};
  gpu_interface_alloc_available_i = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  gpu_interface_cu_id_i = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  gpu_interface_dealloc_wg_id_i = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  dispatch2cu_wf_dispatch_handlers_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dispatch2cu_wf_dispatch_handlers_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  invalid_due_to_not_ready_handlers_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  invalid_due_to_not_ready_handlers_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dispatch2cu_wf_tag_dispatch_handlers_0 = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  dispatch2cu_wf_tag_dispatch_handlers_1 = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  handler_wg_alloc_en_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  handler_wg_alloc_en_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  handler_wg_alloc_wg_id_0 = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  handler_wg_alloc_wg_id_1 = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  handler_wg_alloc_wf_count_0 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  handler_wg_alloc_wf_count_1 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  dispatch2cu_wf_dispatch_i = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  dispatch2cu_wg_wf_count_i = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  dispatch2cu_wf_size_dispatch_i = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  dispatch2cu_sgpr_base_dispatch_i = _RAND_45[12:0];
  _RAND_46 = {1{`RANDOM}};
  dispatch2cu_vgpr_base_dispatch_i = _RAND_46[12:0];
  _RAND_47 = {1{`RANDOM}};
  dispatch2cu_wf_tag_dispatch_i = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  dispatch2cu_lds_base_dispatch_i = _RAND_48[12:0];
  _RAND_49 = {1{`RANDOM}};
  dispatch2cu_start_pc_dispatch_i = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  alloc_st = _RAND_50[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dis_controller(
  input        clock,
  input        reset,
  output       io_dis_controller_start_alloc,
  output       io_dis_controller_alloc_ack,
  output       io_dis_controller_wg_alloc_valid,
  output       io_dis_controller_wg_dealloc_valid,
  output       io_dis_controller_wg_rejected_valid,
  output [1:0] io_dis_controller_cu_busy,
  input        io_inflight_wg_buffer_alloc_valid,
  input        io_inflight_wg_buffer_alloc_available,
  input        io_allocator_cu_valid,
  input        io_allocator_cu_rejected,
  input  [1:0] io_allocator_cu_id_out,
  input        io_grt_wg_alloc_done,
  input        io_grt_wg_dealloc_done,
  input  [1:0] io_grt_wg_alloc_cu_id,
  input  [1:0] io_grt_wg_dealloc_cu_id,
  input        io_gpu_interface_alloc_available,
  input        io_gpu_interface_dealloc_available,
  input  [1:0] io_gpu_interface_cu_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] alloc_st; // @[dis_controller.scala 38:27]
  reg  cu_groups_allocating_0; // @[dis_controller.scala 40:39]
  reg  cu_groups_allocating_1; // @[dis_controller.scala 40:39]
  reg [1:0] alloc_waiting_cu_id; // @[dis_controller.scala 41:38]
  reg  alloc_waiting; // @[dis_controller.scala 42:32]
  reg  dis_controller_start_alloc_i; // @[dis_controller.scala 43:47]
  reg  dis_controller_alloc_ack_i; // @[dis_controller.scala 44:45]
  reg  dis_controller_wg_alloc_valid_i; // @[dis_controller.scala 45:50]
  reg  dis_controller_wg_dealloc_valid_i; // @[dis_controller.scala 46:52]
  reg  dis_controller_wg_rejected_valid_i; // @[dis_controller.scala 47:53]
  wire  gpu_interface_cu_res_tbl_addr = io_gpu_interface_cu_id[1]; // @[dis_controller.scala 54:60]
  wire  _T_5 = io_inflight_wg_buffer_alloc_valid & (~cu_groups_allocating_0 | ~cu_groups_allocating_1); // @[dis_controller.scala 63:52]
  wire  _GEN_2 = io_allocator_cu_valid | alloc_waiting; // @[dis_controller.scala 69:40 70:31 42:32]
  wire  _T_8 = ~alloc_waiting; // @[dis_controller.scala 76:18]
  wire [3:0] _GEN_6 = ~alloc_waiting ? 4'h8 : alloc_st; // @[dis_controller.scala 76:33 78:26 38:27]
  wire [3:0] _GEN_7 = 4'h8 == alloc_st ? 4'h0 : alloc_st; // @[dis_controller.scala 61:21 82:22 38:27]
  wire  _GEN_10 = 4'h2 == alloc_st ? _GEN_2 : alloc_waiting; // @[dis_controller.scala 61:21 42:32]
  wire  _GEN_14 = 4'h0 == alloc_st & _T_5; // @[dis_controller.scala 61:21 57:34]
  wire  _GEN_16 = 4'h0 == alloc_st ? alloc_waiting : _GEN_10; // @[dis_controller.scala 61:21 42:32]
  wire  _GEN_20 = gpu_interface_cu_res_tbl_addr ? cu_groups_allocating_1 : cu_groups_allocating_0; // @[dis_controller.scala 91:{48,48}]
  wire  _T_11 = io_gpu_interface_dealloc_available & ~_GEN_20; // @[dis_controller.scala 91:45]
  wire  _GEN_21 = ~gpu_interface_cu_res_tbl_addr | cu_groups_allocating_0; // @[dis_controller.scala 40:39 93:{61,61}]
  wire  _GEN_22 = gpu_interface_cu_res_tbl_addr | cu_groups_allocating_1; // @[dis_controller.scala 40:39 93:{61,61}]
  wire  _GEN_24 = alloc_waiting_cu_id[1] ? cu_groups_allocating_1 : cu_groups_allocating_0; // @[dis_controller.scala 95:{32,32}]
  wire  _T_15 = io_gpu_interface_alloc_available & io_inflight_wg_buffer_alloc_available; // @[dis_controller.scala 100:52]
  wire  _GEN_25 = ~alloc_waiting_cu_id[1] | cu_groups_allocating_0; // @[dis_controller.scala 103:{108,108} 40:39]
  wire  _GEN_26 = alloc_waiting_cu_id[1] | cu_groups_allocating_1; // @[dis_controller.scala 103:{108,108} 40:39]
  wire  _GEN_27 = io_gpu_interface_alloc_available & io_inflight_wg_buffer_alloc_available ? 1'h0 : _GEN_16; // @[dis_controller.scala 100:93 101:27]
  wire  _GEN_29 = io_gpu_interface_alloc_available & io_inflight_wg_buffer_alloc_available ? _GEN_25 :
    cu_groups_allocating_0; // @[dis_controller.scala 100:93 40:39]
  wire  _GEN_30 = io_gpu_interface_alloc_available & io_inflight_wg_buffer_alloc_available ? _GEN_26 :
    cu_groups_allocating_1; // @[dis_controller.scala 100:93 40:39]
  wire  _GEN_33 = io_allocator_cu_rejected ? 1'h0 : _T_15; // @[dis_controller.scala 96:39 89:41]
  wire  _GEN_34 = io_allocator_cu_rejected ? cu_groups_allocating_0 : _GEN_29; // @[dis_controller.scala 40:39 96:39]
  wire  _GEN_35 = io_allocator_cu_rejected ? cu_groups_allocating_1 : _GEN_30; // @[dis_controller.scala 40:39 96:39]
  wire  _GEN_37 = alloc_waiting & ~_GEN_24 & io_allocator_cu_rejected; // @[dis_controller.scala 95:128 90:44]
  wire  _GEN_38 = alloc_waiting & ~_GEN_24 & _GEN_33; // @[dis_controller.scala 95:128 89:41]
  wire  _GEN_39 = alloc_waiting & ~_GEN_24 ? _GEN_34 : cu_groups_allocating_0; // @[dis_controller.scala 95:128 40:39]
  wire  _GEN_40 = alloc_waiting & ~_GEN_24 ? _GEN_35 : cu_groups_allocating_1; // @[dis_controller.scala 95:128 40:39]
  wire  _GEN_42 = io_gpu_interface_dealloc_available & ~_GEN_20 ? _GEN_21 : _GEN_39; // @[dis_controller.scala 91:101]
  wire  _GEN_43 = io_gpu_interface_dealloc_available & ~_GEN_20 ? _GEN_22 : _GEN_40; // @[dis_controller.scala 91:101]
  assign io_dis_controller_start_alloc = dis_controller_start_alloc_i; // @[dis_controller.scala 48:35]
  assign io_dis_controller_alloc_ack = dis_controller_alloc_ack_i; // @[dis_controller.scala 49:33]
  assign io_dis_controller_wg_alloc_valid = dis_controller_wg_alloc_valid_i; // @[dis_controller.scala 50:38]
  assign io_dis_controller_wg_dealloc_valid = dis_controller_wg_dealloc_valid_i; // @[dis_controller.scala 51:40]
  assign io_dis_controller_wg_rejected_valid = dis_controller_wg_rejected_valid_i; // @[dis_controller.scala 52:41]
  assign io_dis_controller_cu_busy = {cu_groups_allocating_0,cu_groups_allocating_0}; // @[dis_controller.scala 117:49]
  always @(posedge clock) begin
    if (reset) begin // @[dis_controller.scala 38:27]
      alloc_st <= 4'h0; // @[dis_controller.scala 38:27]
    end else if (4'h0 == alloc_st) begin // @[dis_controller.scala 61:21]
      if (io_inflight_wg_buffer_alloc_valid & (~cu_groups_allocating_0 | ~cu_groups_allocating_1)) begin // @[dis_controller.scala 63:94]
        alloc_st <= 4'h2; // @[dis_controller.scala 65:26]
      end
    end else if (4'h2 == alloc_st) begin // @[dis_controller.scala 61:21]
      if (io_allocator_cu_valid) begin // @[dis_controller.scala 69:40]
        alloc_st <= 4'h4; // @[dis_controller.scala 72:26]
      end
    end else if (4'h4 == alloc_st) begin // @[dis_controller.scala 61:21]
      alloc_st <= _GEN_6;
    end else begin
      alloc_st <= _GEN_7;
    end
    if (reset) begin // @[dis_controller.scala 40:39]
      cu_groups_allocating_0 <= 1'h0; // @[dis_controller.scala 40:39]
    end else if (io_grt_wg_alloc_done) begin // @[dis_controller.scala 107:31]
      if (~io_grt_wg_alloc_cu_id[1]) begin // @[dis_controller.scala 108:106]
        cu_groups_allocating_0 <= 1'h0; // @[dis_controller.scala 108:106]
      end else begin
        cu_groups_allocating_0 <= _GEN_42;
      end
    end else if (io_grt_wg_dealloc_done) begin // @[dis_controller.scala 110:38]
      if (~io_grt_wg_dealloc_cu_id[1]) begin // @[dis_controller.scala 111:108]
        cu_groups_allocating_0 <= 1'h0; // @[dis_controller.scala 111:108]
      end else begin
        cu_groups_allocating_0 <= _GEN_42;
      end
    end else begin
      cu_groups_allocating_0 <= _GEN_42;
    end
    if (reset) begin // @[dis_controller.scala 40:39]
      cu_groups_allocating_1 <= 1'h0; // @[dis_controller.scala 40:39]
    end else if (io_grt_wg_alloc_done) begin // @[dis_controller.scala 107:31]
      if (io_grt_wg_alloc_cu_id[1]) begin // @[dis_controller.scala 108:106]
        cu_groups_allocating_1 <= 1'h0; // @[dis_controller.scala 108:106]
      end else begin
        cu_groups_allocating_1 <= _GEN_43;
      end
    end else if (io_grt_wg_dealloc_done) begin // @[dis_controller.scala 110:38]
      if (io_grt_wg_dealloc_cu_id[1]) begin // @[dis_controller.scala 111:108]
        cu_groups_allocating_1 <= 1'h0; // @[dis_controller.scala 111:108]
      end else begin
        cu_groups_allocating_1 <= _GEN_43;
      end
    end else begin
      cu_groups_allocating_1 <= _GEN_43;
    end
    if (reset) begin // @[dis_controller.scala 41:38]
      alloc_waiting_cu_id <= 2'h0; // @[dis_controller.scala 41:38]
    end else if (!(4'h0 == alloc_st)) begin // @[dis_controller.scala 61:21]
      if (4'h2 == alloc_st) begin // @[dis_controller.scala 61:21]
        if (io_allocator_cu_valid) begin // @[dis_controller.scala 69:40]
          alloc_waiting_cu_id <= io_allocator_cu_id_out; // @[dis_controller.scala 71:37]
        end
      end
    end
    if (reset) begin // @[dis_controller.scala 42:32]
      alloc_waiting <= 1'h0; // @[dis_controller.scala 42:32]
    end else if (io_gpu_interface_dealloc_available & ~_GEN_20) begin // @[dis_controller.scala 91:101]
      alloc_waiting <= _GEN_16;
    end else if (alloc_waiting & ~_GEN_24) begin // @[dis_controller.scala 95:128]
      if (io_allocator_cu_rejected) begin // @[dis_controller.scala 96:39]
        alloc_waiting <= 1'h0; // @[dis_controller.scala 97:27]
      end else begin
        alloc_waiting <= _GEN_27;
      end
    end else begin
      alloc_waiting <= _GEN_16;
    end
    if (reset) begin // @[dis_controller.scala 43:47]
      dis_controller_start_alloc_i <= 1'h0; // @[dis_controller.scala 43:47]
    end else begin
      dis_controller_start_alloc_i <= _GEN_14;
    end
    if (reset) begin // @[dis_controller.scala 44:45]
      dis_controller_alloc_ack_i <= 1'h0; // @[dis_controller.scala 44:45]
    end else if (4'h0 == alloc_st) begin // @[dis_controller.scala 61:21]
      dis_controller_alloc_ack_i <= 1'h0; // @[dis_controller.scala 58:32]
    end else if (4'h2 == alloc_st) begin // @[dis_controller.scala 61:21]
      dis_controller_alloc_ack_i <= 1'h0; // @[dis_controller.scala 58:32]
    end else begin
      dis_controller_alloc_ack_i <= 4'h4 == alloc_st & _T_8;
    end
    if (reset) begin // @[dis_controller.scala 45:50]
      dis_controller_wg_alloc_valid_i <= 1'h0; // @[dis_controller.scala 45:50]
    end else if (io_gpu_interface_dealloc_available & ~_GEN_20) begin // @[dis_controller.scala 91:101]
      dis_controller_wg_alloc_valid_i <= 1'h0; // @[dis_controller.scala 89:41]
    end else begin
      dis_controller_wg_alloc_valid_i <= _GEN_38;
    end
    if (reset) begin // @[dis_controller.scala 46:52]
      dis_controller_wg_dealloc_valid_i <= 1'h0; // @[dis_controller.scala 46:52]
    end else begin
      dis_controller_wg_dealloc_valid_i <= _T_11;
    end
    if (reset) begin // @[dis_controller.scala 47:53]
      dis_controller_wg_rejected_valid_i <= 1'h0; // @[dis_controller.scala 47:53]
    end else if (io_gpu_interface_dealloc_available & ~_GEN_20) begin // @[dis_controller.scala 91:101]
      dis_controller_wg_rejected_valid_i <= 1'h0; // @[dis_controller.scala 90:44]
    end else begin
      dis_controller_wg_rejected_valid_i <= _GEN_37;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  alloc_st = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  cu_groups_allocating_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cu_groups_allocating_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alloc_waiting_cu_id = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  alloc_waiting = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dis_controller_start_alloc_i = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dis_controller_alloc_ack_i = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dis_controller_wg_alloc_valid_i = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dis_controller_wg_dealloc_valid_i = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dis_controller_wg_rejected_valid_i = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cta_scheduler(
  input         clock,
  input         reset,
  input         io_host_wg_valid,
  input  [4:0]  io_host_wg_id,
  input  [2:0]  io_host_num_wf,
  input  [9:0]  io_host_wf_size,
  input  [31:0] io_host_start_pc,
  input  [12:0] io_host_vgpr_size_total,
  input  [12:0] io_host_sgpr_size_total,
  input  [12:0] io_host_lds_size_total,
  input  [10:0] io_host_gds_size_total,
  input  [12:0] io_host_vgpr_size_per_wf,
  input  [12:0] io_host_sgpr_size_per_wf,
  output        io_inflight_wg_buffer_host_rcvd_ack,
  output        io_inflight_wg_buffer_host_wf_done,
  output [4:0]  io_inflight_wg_buffer_host_wf_done_wg_id,
  output [1:0]  io_dispatch2cu_wf_dispatch,
  output [2:0]  io_dispatch2cu_wg_wf_count,
  output [9:0]  io_dispatch2cu_wf_size_dispatch,
  output [12:0] io_dispatch2cu_sgpr_base_dispatch,
  output [12:0] io_dispatch2cu_vgpr_base_dispatch,
  output [4:0]  io_dispatch2cu_wf_tag_dispatch,
  output [12:0] io_dispatch2cu_lds_base_dispatch,
  output [31:0] io_dispatch2cu_start_pc_dispatch,
  input  [1:0]  io_cu2dispatch_wf_done,
  input  [4:0]  io_cu2dispatch_wf_tag_done_0,
  input  [4:0]  io_cu2dispatch_wf_tag_done_1,
  input         io_cu2dispatch_ready_for_dispatch_0,
  input         io_cu2dispatch_ready_for_dispatch_1
);
  wire  allocator_neo_i_clock; // @[cta_scheduler.scala 84:33]
  wire  allocator_neo_i_reset; // @[cta_scheduler.scala 84:33]
  wire  allocator_neo_i_io_allocator_cu_valid; // @[cta_scheduler.scala 84:33]
  wire  allocator_neo_i_io_allocator_cu_rejected; // @[cta_scheduler.scala 84:33]
  wire [4:0] allocator_neo_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 84:33]
  wire [1:0] allocator_neo_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 84:33]
  wire [2:0] allocator_neo_i_io_allocator_wf_count; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_allocator_vgpr_size_out; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_allocator_sgpr_size_out; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_allocator_lds_size_out; // @[cta_scheduler.scala 84:33]
  wire [11:0] allocator_neo_i_io_allocator_vgpr_start_out; // @[cta_scheduler.scala 84:33]
  wire [11:0] allocator_neo_i_io_allocator_sgpr_start_out; // @[cta_scheduler.scala 84:33]
  wire [11:0] allocator_neo_i_io_allocator_lds_start_out; // @[cta_scheduler.scala 84:33]
  wire [4:0] allocator_neo_i_io_inflight_wg_buffer_alloc_wg_id; // @[cta_scheduler.scala 84:33]
  wire [2:0] allocator_neo_i_io_inflight_wg_buffer_alloc_num_wf; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_inflight_wg_buffer_alloc_vgpr_size; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_inflight_wg_buffer_alloc_sgpr_size; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_inflight_wg_buffer_alloc_lds_size; // @[cta_scheduler.scala 84:33]
  wire [1:0] allocator_neo_i_io_dis_controller_cu_busy; // @[cta_scheduler.scala 84:33]
  wire  allocator_neo_i_io_dis_controller_alloc_ack; // @[cta_scheduler.scala 84:33]
  wire  allocator_neo_i_io_dis_controller_start_alloc; // @[cta_scheduler.scala 84:33]
  wire  allocator_neo_i_io_grt_cam_up_valid; // @[cta_scheduler.scala 84:33]
  wire [1:0] allocator_neo_i_io_grt_cam_up_cu_id; // @[cta_scheduler.scala 84:33]
  wire [11:0] allocator_neo_i_io_grt_cam_up_vgpr_strt; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_grt_cam_up_vgpr_size; // @[cta_scheduler.scala 84:33]
  wire [11:0] allocator_neo_i_io_grt_cam_up_sgpr_strt; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_grt_cam_up_sgpr_size; // @[cta_scheduler.scala 84:33]
  wire [11:0] allocator_neo_i_io_grt_cam_up_lds_strt; // @[cta_scheduler.scala 84:33]
  wire [12:0] allocator_neo_i_io_grt_cam_up_lds_size; // @[cta_scheduler.scala 84:33]
  wire [2:0] allocator_neo_i_io_grt_cam_up_wf_count; // @[cta_scheduler.scala 84:33]
  wire [2:0] allocator_neo_i_io_grt_cam_up_wg_count; // @[cta_scheduler.scala 84:33]
  wire  top_resource_table_i_clock; // @[cta_scheduler.scala 85:38]
  wire  top_resource_table_i_reset; // @[cta_scheduler.scala 85:38]
  wire  top_resource_table_i_io_grt_cam_up_valid; // @[cta_scheduler.scala 85:38]
  wire [2:0] top_resource_table_i_io_grt_cam_up_wf_count; // @[cta_scheduler.scala 85:38]
  wire [1:0] top_resource_table_i_io_grt_cam_up_cu_id; // @[cta_scheduler.scala 85:38]
  wire [11:0] top_resource_table_i_io_grt_cam_up_vgpr_strt; // @[cta_scheduler.scala 85:38]
  wire [12:0] top_resource_table_i_io_grt_cam_up_vgpr_size; // @[cta_scheduler.scala 85:38]
  wire [11:0] top_resource_table_i_io_grt_cam_up_sgpr_strt; // @[cta_scheduler.scala 85:38]
  wire [12:0] top_resource_table_i_io_grt_cam_up_sgpr_size; // @[cta_scheduler.scala 85:38]
  wire [11:0] top_resource_table_i_io_grt_cam_up_lds_strt; // @[cta_scheduler.scala 85:38]
  wire [12:0] top_resource_table_i_io_grt_cam_up_lds_size; // @[cta_scheduler.scala 85:38]
  wire [2:0] top_resource_table_i_io_grt_cam_up_wg_count; // @[cta_scheduler.scala 85:38]
  wire  top_resource_table_i_io_grt_wg_alloc_done; // @[cta_scheduler.scala 85:38]
  wire [1:0] top_resource_table_i_io_grt_wg_alloc_cu_id; // @[cta_scheduler.scala 85:38]
  wire  top_resource_table_i_io_grt_wg_dealloc_done; // @[cta_scheduler.scala 85:38]
  wire [1:0] top_resource_table_i_io_grt_wg_dealloc_cu_id; // @[cta_scheduler.scala 85:38]
  wire [1:0] top_resource_table_i_io_gpu_interface_cu_id; // @[cta_scheduler.scala 85:38]
  wire [4:0] top_resource_table_i_io_gpu_interface_dealloc_wg_id; // @[cta_scheduler.scala 85:38]
  wire  top_resource_table_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 85:38]
  wire  top_resource_table_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 85:38]
  wire [4:0] top_resource_table_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 85:38]
  wire [2:0] top_resource_table_i_io_allocator_wf_count; // @[cta_scheduler.scala 85:38]
  wire [1:0] top_resource_table_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 85:38]
  wire [11:0] top_resource_table_i_io_allocator_vgpr_start_out; // @[cta_scheduler.scala 85:38]
  wire [12:0] top_resource_table_i_io_allocator_vgpr_size_out; // @[cta_scheduler.scala 85:38]
  wire [11:0] top_resource_table_i_io_allocator_sgpr_start_out; // @[cta_scheduler.scala 85:38]
  wire [12:0] top_resource_table_i_io_allocator_sgpr_size_out; // @[cta_scheduler.scala 85:38]
  wire [11:0] top_resource_table_i_io_allocator_lds_start_out; // @[cta_scheduler.scala 85:38]
  wire [12:0] top_resource_table_i_io_allocator_lds_size_out; // @[cta_scheduler.scala 85:38]
  wire  inflight_wg_buffer_i_clock; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_reset; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_host_wg_valid; // @[cta_scheduler.scala 86:38]
  wire [4:0] inflight_wg_buffer_i_io_host_wg_id; // @[cta_scheduler.scala 86:38]
  wire [2:0] inflight_wg_buffer_i_io_host_num_wf; // @[cta_scheduler.scala 86:38]
  wire [9:0] inflight_wg_buffer_i_io_host_wf_size; // @[cta_scheduler.scala 86:38]
  wire [31:0] inflight_wg_buffer_i_io_host_start_pc; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_host_vgpr_size_total; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_host_sgpr_size_total; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_host_lds_size_total; // @[cta_scheduler.scala 86:38]
  wire [10:0] inflight_wg_buffer_i_io_host_gds_size_total; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_host_vgpr_size_per_wf; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_host_sgpr_size_per_wf; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_dis_controller_start_alloc; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_dis_controller_wg_rejected_valid; // @[cta_scheduler.scala 86:38]
  wire [4:0] inflight_wg_buffer_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 86:38]
  wire [4:0] inflight_wg_buffer_i_io_gpu_interface_dealloc_wg_id; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_inflight_wg_buffer_host_rcvd_ack; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_inflight_wg_buffer_host_wf_done; // @[cta_scheduler.scala 86:38]
  wire [4:0] inflight_wg_buffer_i_io_inflight_wg_buffer_host_wf_done_wg_id; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_valid; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_available; // @[cta_scheduler.scala 86:38]
  wire [4:0] inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_wg_id; // @[cta_scheduler.scala 86:38]
  wire [2:0] inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_num_wf; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_vgpr_size; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_sgpr_size; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_lds_size; // @[cta_scheduler.scala 86:38]
  wire  inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_valid; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_vgpr_size_per_wf; // @[cta_scheduler.scala 86:38]
  wire [12:0] inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_sgpr_size_per_wf; // @[cta_scheduler.scala 86:38]
  wire [9:0] inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_wf_size; // @[cta_scheduler.scala 86:38]
  wire [31:0] inflight_wg_buffer_i_io_inflight_wg_buffer_start_pc; // @[cta_scheduler.scala 86:38]
  wire  gpu_interface_i_clock; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_reset; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_inflight_wg_buffer_gpu_valid; // @[cta_scheduler.scala 87:33]
  wire [9:0] gpu_interface_i_io_inflight_wg_buffer_gpu_wf_size; // @[cta_scheduler.scala 87:33]
  wire [31:0] gpu_interface_i_io_inflight_wg_buffer_start_pc; // @[cta_scheduler.scala 87:33]
  wire [11:0] gpu_interface_i_io_inflight_wg_buffer_gpu_vgpr_size_per_wf; // @[cta_scheduler.scala 87:33]
  wire [11:0] gpu_interface_i_io_inflight_wg_buffer_gpu_sgpr_size_per_wf; // @[cta_scheduler.scala 87:33]
  wire [4:0] gpu_interface_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 87:33]
  wire [1:0] gpu_interface_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 87:33]
  wire [2:0] gpu_interface_i_io_allocator_wf_count; // @[cta_scheduler.scala 87:33]
  wire [11:0] gpu_interface_i_io_allocator_vgpr_start_out; // @[cta_scheduler.scala 87:33]
  wire [11:0] gpu_interface_i_io_allocator_sgpr_start_out; // @[cta_scheduler.scala 87:33]
  wire [11:0] gpu_interface_i_io_allocator_lds_start_out; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_gpu_interface_alloc_available; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_gpu_interface_dealloc_available; // @[cta_scheduler.scala 87:33]
  wire [1:0] gpu_interface_i_io_gpu_interface_cu_id; // @[cta_scheduler.scala 87:33]
  wire [4:0] gpu_interface_i_io_gpu_interface_dealloc_wg_id; // @[cta_scheduler.scala 87:33]
  wire [1:0] gpu_interface_i_io_dispatch2cu_wf_dispatch; // @[cta_scheduler.scala 87:33]
  wire [2:0] gpu_interface_i_io_dispatch2cu_wg_wf_count; // @[cta_scheduler.scala 87:33]
  wire [9:0] gpu_interface_i_io_dispatch2cu_wf_size_dispatch; // @[cta_scheduler.scala 87:33]
  wire [12:0] gpu_interface_i_io_dispatch2cu_sgpr_base_dispatch; // @[cta_scheduler.scala 87:33]
  wire [12:0] gpu_interface_i_io_dispatch2cu_vgpr_base_dispatch; // @[cta_scheduler.scala 87:33]
  wire [4:0] gpu_interface_i_io_dispatch2cu_wf_tag_dispatch; // @[cta_scheduler.scala 87:33]
  wire [12:0] gpu_interface_i_io_dispatch2cu_lds_base_dispatch; // @[cta_scheduler.scala 87:33]
  wire [31:0] gpu_interface_i_io_dispatch2cu_start_pc_dispatch; // @[cta_scheduler.scala 87:33]
  wire [1:0] gpu_interface_i_io_cu2dispatch_wf_done; // @[cta_scheduler.scala 87:33]
  wire [4:0] gpu_interface_i_io_cu2dispatch_wf_tag_done_0; // @[cta_scheduler.scala 87:33]
  wire [4:0] gpu_interface_i_io_cu2dispatch_wf_tag_done_1; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_cu2dispatch_ready_for_dispatch_0; // @[cta_scheduler.scala 87:33]
  wire  gpu_interface_i_io_cu2dispatch_ready_for_dispatch_1; // @[cta_scheduler.scala 87:33]
  wire  dis_controller_i_clock; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_reset; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_dis_controller_start_alloc; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_dis_controller_alloc_ack; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_dis_controller_wg_rejected_valid; // @[cta_scheduler.scala 88:34]
  wire [1:0] dis_controller_i_io_dis_controller_cu_busy; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_inflight_wg_buffer_alloc_valid; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_inflight_wg_buffer_alloc_available; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_allocator_cu_valid; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_allocator_cu_rejected; // @[cta_scheduler.scala 88:34]
  wire [1:0] dis_controller_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_grt_wg_alloc_done; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_grt_wg_dealloc_done; // @[cta_scheduler.scala 88:34]
  wire [1:0] dis_controller_i_io_grt_wg_alloc_cu_id; // @[cta_scheduler.scala 88:34]
  wire [1:0] dis_controller_i_io_grt_wg_dealloc_cu_id; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_gpu_interface_alloc_available; // @[cta_scheduler.scala 88:34]
  wire  dis_controller_i_io_gpu_interface_dealloc_available; // @[cta_scheduler.scala 88:34]
  wire [1:0] dis_controller_i_io_gpu_interface_cu_id; // @[cta_scheduler.scala 88:34]
  wire [12:0] inflight_wg_buffer_gpu_vgpr_size_per_wf = inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_vgpr_size_per_wf; // @[cta_scheduler.scala 146:45 48:55]
  wire [12:0] inflight_wg_buffer_gpu_sgpr_size_per_wf = inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_sgpr_size_per_wf; // @[cta_scheduler.scala 147:45 49:55]
  wire [11:0] allocator_vgpr_size_out = allocator_neo_i_io_allocator_vgpr_size_out[11:0]; // @[cta_scheduler.scala 76:39 94:29]
  wire [11:0] allocator_sgpr_size_out = allocator_neo_i_io_allocator_sgpr_size_out[11:0]; // @[cta_scheduler.scala 77:39 95:29]
  wire [11:0] allocator_lds_size_out = allocator_neo_i_io_allocator_lds_size_out[11:0]; // @[cta_scheduler.scala 78:38 96:28]
  allocator_neo allocator_neo_i ( // @[cta_scheduler.scala 84:33]
    .clock(allocator_neo_i_clock),
    .reset(allocator_neo_i_reset),
    .io_allocator_cu_valid(allocator_neo_i_io_allocator_cu_valid),
    .io_allocator_cu_rejected(allocator_neo_i_io_allocator_cu_rejected),
    .io_allocator_wg_id_out(allocator_neo_i_io_allocator_wg_id_out),
    .io_allocator_cu_id_out(allocator_neo_i_io_allocator_cu_id_out),
    .io_allocator_wf_count(allocator_neo_i_io_allocator_wf_count),
    .io_allocator_vgpr_size_out(allocator_neo_i_io_allocator_vgpr_size_out),
    .io_allocator_sgpr_size_out(allocator_neo_i_io_allocator_sgpr_size_out),
    .io_allocator_lds_size_out(allocator_neo_i_io_allocator_lds_size_out),
    .io_allocator_vgpr_start_out(allocator_neo_i_io_allocator_vgpr_start_out),
    .io_allocator_sgpr_start_out(allocator_neo_i_io_allocator_sgpr_start_out),
    .io_allocator_lds_start_out(allocator_neo_i_io_allocator_lds_start_out),
    .io_inflight_wg_buffer_alloc_wg_id(allocator_neo_i_io_inflight_wg_buffer_alloc_wg_id),
    .io_inflight_wg_buffer_alloc_num_wf(allocator_neo_i_io_inflight_wg_buffer_alloc_num_wf),
    .io_inflight_wg_buffer_alloc_vgpr_size(allocator_neo_i_io_inflight_wg_buffer_alloc_vgpr_size),
    .io_inflight_wg_buffer_alloc_sgpr_size(allocator_neo_i_io_inflight_wg_buffer_alloc_sgpr_size),
    .io_inflight_wg_buffer_alloc_lds_size(allocator_neo_i_io_inflight_wg_buffer_alloc_lds_size),
    .io_dis_controller_cu_busy(allocator_neo_i_io_dis_controller_cu_busy),
    .io_dis_controller_alloc_ack(allocator_neo_i_io_dis_controller_alloc_ack),
    .io_dis_controller_start_alloc(allocator_neo_i_io_dis_controller_start_alloc),
    .io_grt_cam_up_valid(allocator_neo_i_io_grt_cam_up_valid),
    .io_grt_cam_up_cu_id(allocator_neo_i_io_grt_cam_up_cu_id),
    .io_grt_cam_up_vgpr_strt(allocator_neo_i_io_grt_cam_up_vgpr_strt),
    .io_grt_cam_up_vgpr_size(allocator_neo_i_io_grt_cam_up_vgpr_size),
    .io_grt_cam_up_sgpr_strt(allocator_neo_i_io_grt_cam_up_sgpr_strt),
    .io_grt_cam_up_sgpr_size(allocator_neo_i_io_grt_cam_up_sgpr_size),
    .io_grt_cam_up_lds_strt(allocator_neo_i_io_grt_cam_up_lds_strt),
    .io_grt_cam_up_lds_size(allocator_neo_i_io_grt_cam_up_lds_size),
    .io_grt_cam_up_wf_count(allocator_neo_i_io_grt_cam_up_wf_count),
    .io_grt_cam_up_wg_count(allocator_neo_i_io_grt_cam_up_wg_count)
  );
  top_resource_table top_resource_table_i ( // @[cta_scheduler.scala 85:38]
    .clock(top_resource_table_i_clock),
    .reset(top_resource_table_i_reset),
    .io_grt_cam_up_valid(top_resource_table_i_io_grt_cam_up_valid),
    .io_grt_cam_up_wf_count(top_resource_table_i_io_grt_cam_up_wf_count),
    .io_grt_cam_up_cu_id(top_resource_table_i_io_grt_cam_up_cu_id),
    .io_grt_cam_up_vgpr_strt(top_resource_table_i_io_grt_cam_up_vgpr_strt),
    .io_grt_cam_up_vgpr_size(top_resource_table_i_io_grt_cam_up_vgpr_size),
    .io_grt_cam_up_sgpr_strt(top_resource_table_i_io_grt_cam_up_sgpr_strt),
    .io_grt_cam_up_sgpr_size(top_resource_table_i_io_grt_cam_up_sgpr_size),
    .io_grt_cam_up_lds_strt(top_resource_table_i_io_grt_cam_up_lds_strt),
    .io_grt_cam_up_lds_size(top_resource_table_i_io_grt_cam_up_lds_size),
    .io_grt_cam_up_wg_count(top_resource_table_i_io_grt_cam_up_wg_count),
    .io_grt_wg_alloc_done(top_resource_table_i_io_grt_wg_alloc_done),
    .io_grt_wg_alloc_cu_id(top_resource_table_i_io_grt_wg_alloc_cu_id),
    .io_grt_wg_dealloc_done(top_resource_table_i_io_grt_wg_dealloc_done),
    .io_grt_wg_dealloc_cu_id(top_resource_table_i_io_grt_wg_dealloc_cu_id),
    .io_gpu_interface_cu_id(top_resource_table_i_io_gpu_interface_cu_id),
    .io_gpu_interface_dealloc_wg_id(top_resource_table_i_io_gpu_interface_dealloc_wg_id),
    .io_dis_controller_wg_alloc_valid(top_resource_table_i_io_dis_controller_wg_alloc_valid),
    .io_dis_controller_wg_dealloc_valid(top_resource_table_i_io_dis_controller_wg_dealloc_valid),
    .io_allocator_wg_id_out(top_resource_table_i_io_allocator_wg_id_out),
    .io_allocator_wf_count(top_resource_table_i_io_allocator_wf_count),
    .io_allocator_cu_id_out(top_resource_table_i_io_allocator_cu_id_out),
    .io_allocator_vgpr_start_out(top_resource_table_i_io_allocator_vgpr_start_out),
    .io_allocator_vgpr_size_out(top_resource_table_i_io_allocator_vgpr_size_out),
    .io_allocator_sgpr_start_out(top_resource_table_i_io_allocator_sgpr_start_out),
    .io_allocator_sgpr_size_out(top_resource_table_i_io_allocator_sgpr_size_out),
    .io_allocator_lds_start_out(top_resource_table_i_io_allocator_lds_start_out),
    .io_allocator_lds_size_out(top_resource_table_i_io_allocator_lds_size_out)
  );
  inflight_wg_buffer inflight_wg_buffer_i ( // @[cta_scheduler.scala 86:38]
    .clock(inflight_wg_buffer_i_clock),
    .reset(inflight_wg_buffer_i_reset),
    .io_host_wg_valid(inflight_wg_buffer_i_io_host_wg_valid),
    .io_host_wg_id(inflight_wg_buffer_i_io_host_wg_id),
    .io_host_num_wf(inflight_wg_buffer_i_io_host_num_wf),
    .io_host_wf_size(inflight_wg_buffer_i_io_host_wf_size),
    .io_host_start_pc(inflight_wg_buffer_i_io_host_start_pc),
    .io_host_vgpr_size_total(inflight_wg_buffer_i_io_host_vgpr_size_total),
    .io_host_sgpr_size_total(inflight_wg_buffer_i_io_host_sgpr_size_total),
    .io_host_lds_size_total(inflight_wg_buffer_i_io_host_lds_size_total),
    .io_host_gds_size_total(inflight_wg_buffer_i_io_host_gds_size_total),
    .io_host_vgpr_size_per_wf(inflight_wg_buffer_i_io_host_vgpr_size_per_wf),
    .io_host_sgpr_size_per_wf(inflight_wg_buffer_i_io_host_sgpr_size_per_wf),
    .io_dis_controller_wg_alloc_valid(inflight_wg_buffer_i_io_dis_controller_wg_alloc_valid),
    .io_dis_controller_start_alloc(inflight_wg_buffer_i_io_dis_controller_start_alloc),
    .io_dis_controller_wg_dealloc_valid(inflight_wg_buffer_i_io_dis_controller_wg_dealloc_valid),
    .io_dis_controller_wg_rejected_valid(inflight_wg_buffer_i_io_dis_controller_wg_rejected_valid),
    .io_allocator_wg_id_out(inflight_wg_buffer_i_io_allocator_wg_id_out),
    .io_gpu_interface_dealloc_wg_id(inflight_wg_buffer_i_io_gpu_interface_dealloc_wg_id),
    .io_inflight_wg_buffer_host_rcvd_ack(inflight_wg_buffer_i_io_inflight_wg_buffer_host_rcvd_ack),
    .io_inflight_wg_buffer_host_wf_done(inflight_wg_buffer_i_io_inflight_wg_buffer_host_wf_done),
    .io_inflight_wg_buffer_host_wf_done_wg_id(inflight_wg_buffer_i_io_inflight_wg_buffer_host_wf_done_wg_id),
    .io_inflight_wg_buffer_alloc_valid(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_valid),
    .io_inflight_wg_buffer_alloc_available(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_available),
    .io_inflight_wg_buffer_alloc_wg_id(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_wg_id),
    .io_inflight_wg_buffer_alloc_num_wf(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_num_wf),
    .io_inflight_wg_buffer_alloc_vgpr_size(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_vgpr_size),
    .io_inflight_wg_buffer_alloc_sgpr_size(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_sgpr_size),
    .io_inflight_wg_buffer_alloc_lds_size(inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_lds_size),
    .io_inflight_wg_buffer_gpu_valid(inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_valid),
    .io_inflight_wg_buffer_gpu_vgpr_size_per_wf(inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_vgpr_size_per_wf),
    .io_inflight_wg_buffer_gpu_sgpr_size_per_wf(inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_sgpr_size_per_wf),
    .io_inflight_wg_buffer_gpu_wf_size(inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_wf_size),
    .io_inflight_wg_buffer_start_pc(inflight_wg_buffer_i_io_inflight_wg_buffer_start_pc)
  );
  gpu_interface gpu_interface_i ( // @[cta_scheduler.scala 87:33]
    .clock(gpu_interface_i_clock),
    .reset(gpu_interface_i_reset),
    .io_inflight_wg_buffer_gpu_valid(gpu_interface_i_io_inflight_wg_buffer_gpu_valid),
    .io_inflight_wg_buffer_gpu_wf_size(gpu_interface_i_io_inflight_wg_buffer_gpu_wf_size),
    .io_inflight_wg_buffer_start_pc(gpu_interface_i_io_inflight_wg_buffer_start_pc),
    .io_inflight_wg_buffer_gpu_vgpr_size_per_wf(gpu_interface_i_io_inflight_wg_buffer_gpu_vgpr_size_per_wf),
    .io_inflight_wg_buffer_gpu_sgpr_size_per_wf(gpu_interface_i_io_inflight_wg_buffer_gpu_sgpr_size_per_wf),
    .io_allocator_wg_id_out(gpu_interface_i_io_allocator_wg_id_out),
    .io_allocator_cu_id_out(gpu_interface_i_io_allocator_cu_id_out),
    .io_allocator_wf_count(gpu_interface_i_io_allocator_wf_count),
    .io_allocator_vgpr_start_out(gpu_interface_i_io_allocator_vgpr_start_out),
    .io_allocator_sgpr_start_out(gpu_interface_i_io_allocator_sgpr_start_out),
    .io_allocator_lds_start_out(gpu_interface_i_io_allocator_lds_start_out),
    .io_dis_controller_wg_alloc_valid(gpu_interface_i_io_dis_controller_wg_alloc_valid),
    .io_dis_controller_wg_dealloc_valid(gpu_interface_i_io_dis_controller_wg_dealloc_valid),
    .io_gpu_interface_alloc_available(gpu_interface_i_io_gpu_interface_alloc_available),
    .io_gpu_interface_dealloc_available(gpu_interface_i_io_gpu_interface_dealloc_available),
    .io_gpu_interface_cu_id(gpu_interface_i_io_gpu_interface_cu_id),
    .io_gpu_interface_dealloc_wg_id(gpu_interface_i_io_gpu_interface_dealloc_wg_id),
    .io_dispatch2cu_wf_dispatch(gpu_interface_i_io_dispatch2cu_wf_dispatch),
    .io_dispatch2cu_wg_wf_count(gpu_interface_i_io_dispatch2cu_wg_wf_count),
    .io_dispatch2cu_wf_size_dispatch(gpu_interface_i_io_dispatch2cu_wf_size_dispatch),
    .io_dispatch2cu_sgpr_base_dispatch(gpu_interface_i_io_dispatch2cu_sgpr_base_dispatch),
    .io_dispatch2cu_vgpr_base_dispatch(gpu_interface_i_io_dispatch2cu_vgpr_base_dispatch),
    .io_dispatch2cu_wf_tag_dispatch(gpu_interface_i_io_dispatch2cu_wf_tag_dispatch),
    .io_dispatch2cu_lds_base_dispatch(gpu_interface_i_io_dispatch2cu_lds_base_dispatch),
    .io_dispatch2cu_start_pc_dispatch(gpu_interface_i_io_dispatch2cu_start_pc_dispatch),
    .io_cu2dispatch_wf_done(gpu_interface_i_io_cu2dispatch_wf_done),
    .io_cu2dispatch_wf_tag_done_0(gpu_interface_i_io_cu2dispatch_wf_tag_done_0),
    .io_cu2dispatch_wf_tag_done_1(gpu_interface_i_io_cu2dispatch_wf_tag_done_1),
    .io_cu2dispatch_ready_for_dispatch_0(gpu_interface_i_io_cu2dispatch_ready_for_dispatch_0),
    .io_cu2dispatch_ready_for_dispatch_1(gpu_interface_i_io_cu2dispatch_ready_for_dispatch_1)
  );
  dis_controller dis_controller_i ( // @[cta_scheduler.scala 88:34]
    .clock(dis_controller_i_clock),
    .reset(dis_controller_i_reset),
    .io_dis_controller_start_alloc(dis_controller_i_io_dis_controller_start_alloc),
    .io_dis_controller_alloc_ack(dis_controller_i_io_dis_controller_alloc_ack),
    .io_dis_controller_wg_alloc_valid(dis_controller_i_io_dis_controller_wg_alloc_valid),
    .io_dis_controller_wg_dealloc_valid(dis_controller_i_io_dis_controller_wg_dealloc_valid),
    .io_dis_controller_wg_rejected_valid(dis_controller_i_io_dis_controller_wg_rejected_valid),
    .io_dis_controller_cu_busy(dis_controller_i_io_dis_controller_cu_busy),
    .io_inflight_wg_buffer_alloc_valid(dis_controller_i_io_inflight_wg_buffer_alloc_valid),
    .io_inflight_wg_buffer_alloc_available(dis_controller_i_io_inflight_wg_buffer_alloc_available),
    .io_allocator_cu_valid(dis_controller_i_io_allocator_cu_valid),
    .io_allocator_cu_rejected(dis_controller_i_io_allocator_cu_rejected),
    .io_allocator_cu_id_out(dis_controller_i_io_allocator_cu_id_out),
    .io_grt_wg_alloc_done(dis_controller_i_io_grt_wg_alloc_done),
    .io_grt_wg_dealloc_done(dis_controller_i_io_grt_wg_dealloc_done),
    .io_grt_wg_alloc_cu_id(dis_controller_i_io_grt_wg_alloc_cu_id),
    .io_grt_wg_dealloc_cu_id(dis_controller_i_io_grt_wg_dealloc_cu_id),
    .io_gpu_interface_alloc_available(dis_controller_i_io_gpu_interface_alloc_available),
    .io_gpu_interface_dealloc_available(dis_controller_i_io_gpu_interface_dealloc_available),
    .io_gpu_interface_cu_id(dis_controller_i_io_gpu_interface_cu_id)
  );
  assign io_inflight_wg_buffer_host_rcvd_ack = inflight_wg_buffer_i_io_inflight_wg_buffer_host_rcvd_ack; // @[cta_scheduler.scala 135:41]
  assign io_inflight_wg_buffer_host_wf_done = inflight_wg_buffer_i_io_inflight_wg_buffer_host_wf_done; // @[cta_scheduler.scala 136:40]
  assign io_inflight_wg_buffer_host_wf_done_wg_id = inflight_wg_buffer_i_io_inflight_wg_buffer_host_wf_done_wg_id; // @[cta_scheduler.scala 137:46]
  assign io_dispatch2cu_wf_dispatch = gpu_interface_i_io_dispatch2cu_wf_dispatch; // @[cta_scheduler.scala 167:32]
  assign io_dispatch2cu_wg_wf_count = gpu_interface_i_io_dispatch2cu_wg_wf_count; // @[cta_scheduler.scala 168:32]
  assign io_dispatch2cu_wf_size_dispatch = gpu_interface_i_io_dispatch2cu_wf_size_dispatch; // @[cta_scheduler.scala 169:37]
  assign io_dispatch2cu_sgpr_base_dispatch = gpu_interface_i_io_dispatch2cu_sgpr_base_dispatch; // @[cta_scheduler.scala 170:39]
  assign io_dispatch2cu_vgpr_base_dispatch = gpu_interface_i_io_dispatch2cu_vgpr_base_dispatch; // @[cta_scheduler.scala 171:39]
  assign io_dispatch2cu_wf_tag_dispatch = gpu_interface_i_io_dispatch2cu_wf_tag_dispatch; // @[cta_scheduler.scala 172:36]
  assign io_dispatch2cu_lds_base_dispatch = gpu_interface_i_io_dispatch2cu_lds_base_dispatch; // @[cta_scheduler.scala 173:38]
  assign io_dispatch2cu_start_pc_dispatch = gpu_interface_i_io_dispatch2cu_start_pc_dispatch; // @[cta_scheduler.scala 174:38]
  assign allocator_neo_i_clock = clock;
  assign allocator_neo_i_reset = reset;
  assign allocator_neo_i_io_inflight_wg_buffer_alloc_wg_id = inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_wg_id; // @[cta_scheduler.scala 140:36 42:46]
  assign allocator_neo_i_io_inflight_wg_buffer_alloc_num_wf = inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_num_wf; // @[cta_scheduler.scala 141:37 43:47]
  assign allocator_neo_i_io_inflight_wg_buffer_alloc_vgpr_size =
    inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_vgpr_size; // @[cta_scheduler.scala 142:40 44:50]
  assign allocator_neo_i_io_inflight_wg_buffer_alloc_sgpr_size =
    inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_sgpr_size; // @[cta_scheduler.scala 143:40 45:50]
  assign allocator_neo_i_io_inflight_wg_buffer_alloc_lds_size =
    inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_lds_size; // @[cta_scheduler.scala 144:39 46:49]
  assign allocator_neo_i_io_dis_controller_cu_busy = dis_controller_i_io_dis_controller_cu_busy; // @[cta_scheduler.scala 212:28 80:38]
  assign allocator_neo_i_io_dis_controller_alloc_ack = dis_controller_i_io_dis_controller_alloc_ack; // @[cta_scheduler.scala 208:30 79:40]
  assign allocator_neo_i_io_dis_controller_start_alloc = dis_controller_i_io_dis_controller_start_alloc; // @[cta_scheduler.scala 207:32 35:42]
  assign allocator_neo_i_io_grt_cam_up_valid = top_resource_table_i_io_grt_cam_up_valid; // @[cta_scheduler.scala 178:22 60:32]
  assign allocator_neo_i_io_grt_cam_up_cu_id = top_resource_table_i_io_grt_cam_up_cu_id; // @[cta_scheduler.scala 181:22 63:32]
  assign allocator_neo_i_io_grt_cam_up_vgpr_strt = top_resource_table_i_io_grt_cam_up_vgpr_strt; // @[cta_scheduler.scala 182:26 64:36]
  assign allocator_neo_i_io_grt_cam_up_vgpr_size = top_resource_table_i_io_grt_cam_up_vgpr_size; // @[cta_scheduler.scala 183:26 65:36]
  assign allocator_neo_i_io_grt_cam_up_sgpr_strt = top_resource_table_i_io_grt_cam_up_sgpr_strt; // @[cta_scheduler.scala 184:26 66:36]
  assign allocator_neo_i_io_grt_cam_up_sgpr_size = top_resource_table_i_io_grt_cam_up_sgpr_size; // @[cta_scheduler.scala 185:26 67:36]
  assign allocator_neo_i_io_grt_cam_up_lds_strt = top_resource_table_i_io_grt_cam_up_lds_strt; // @[cta_scheduler.scala 186:25 68:35]
  assign allocator_neo_i_io_grt_cam_up_lds_size = top_resource_table_i_io_grt_cam_up_lds_size; // @[cta_scheduler.scala 187:25 69:35]
  assign allocator_neo_i_io_grt_cam_up_wf_count = top_resource_table_i_io_grt_cam_up_wf_count; // @[cta_scheduler.scala 179:25 61:35]
  assign allocator_neo_i_io_grt_cam_up_wg_count = top_resource_table_i_io_grt_cam_up_wg_count; // @[cta_scheduler.scala 180:25 62:35]
  assign top_resource_table_i_clock = clock;
  assign top_resource_table_i_reset = reset;
  assign top_resource_table_i_io_gpu_interface_cu_id = gpu_interface_i_io_gpu_interface_cu_id; // @[cta_scheduler.scala 165:25 59:35]
  assign top_resource_table_i_io_gpu_interface_dealloc_wg_id = gpu_interface_i_io_gpu_interface_dealloc_wg_id; // @[cta_scheduler.scala 166:33 39:43]
  assign top_resource_table_i_io_dis_controller_wg_alloc_valid = dis_controller_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 209:35 34:45]
  assign top_resource_table_i_io_dis_controller_wg_dealloc_valid = dis_controller_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 210:37 36:47]
  assign top_resource_table_i_io_allocator_wg_id_out = allocator_neo_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 38:35 91:25]
  assign top_resource_table_i_io_allocator_wf_count = allocator_neo_i_io_allocator_wf_count; // @[cta_scheduler.scala 53:34 93:24]
  assign top_resource_table_i_io_allocator_cu_id_out = allocator_neo_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 52:35 92:25]
  assign top_resource_table_i_io_allocator_vgpr_start_out = allocator_neo_i_io_allocator_vgpr_start_out; // @[cta_scheduler.scala 54:40 97:30]
  assign top_resource_table_i_io_allocator_vgpr_size_out = {{1'd0}, allocator_vgpr_size_out}; // @[cta_scheduler.scala 202:53]
  assign top_resource_table_i_io_allocator_sgpr_start_out = allocator_neo_i_io_allocator_sgpr_start_out; // @[cta_scheduler.scala 55:40 98:30]
  assign top_resource_table_i_io_allocator_sgpr_size_out = {{1'd0}, allocator_sgpr_size_out}; // @[cta_scheduler.scala 204:53]
  assign top_resource_table_i_io_allocator_lds_start_out = allocator_neo_i_io_allocator_lds_start_out; // @[cta_scheduler.scala 56:39 99:29]
  assign top_resource_table_i_io_allocator_lds_size_out = {{1'd0}, allocator_lds_size_out}; // @[cta_scheduler.scala 206:52]
  assign inflight_wg_buffer_i_clock = clock;
  assign inflight_wg_buffer_i_reset = reset;
  assign inflight_wg_buffer_i_io_host_wg_valid = io_host_wg_valid; // @[cta_scheduler.scala 118:43]
  assign inflight_wg_buffer_i_io_host_wg_id = io_host_wg_id; // @[cta_scheduler.scala 119:40]
  assign inflight_wg_buffer_i_io_host_num_wf = io_host_num_wf; // @[cta_scheduler.scala 120:41]
  assign inflight_wg_buffer_i_io_host_wf_size = io_host_wf_size; // @[cta_scheduler.scala 121:42]
  assign inflight_wg_buffer_i_io_host_start_pc = io_host_start_pc; // @[cta_scheduler.scala 122:43]
  assign inflight_wg_buffer_i_io_host_vgpr_size_total = io_host_vgpr_size_total; // @[cta_scheduler.scala 123:50]
  assign inflight_wg_buffer_i_io_host_sgpr_size_total = io_host_sgpr_size_total; // @[cta_scheduler.scala 124:50]
  assign inflight_wg_buffer_i_io_host_lds_size_total = io_host_lds_size_total; // @[cta_scheduler.scala 125:49]
  assign inflight_wg_buffer_i_io_host_gds_size_total = io_host_gds_size_total; // @[cta_scheduler.scala 126:49]
  assign inflight_wg_buffer_i_io_host_vgpr_size_per_wf = io_host_vgpr_size_per_wf; // @[cta_scheduler.scala 127:51]
  assign inflight_wg_buffer_i_io_host_sgpr_size_per_wf = io_host_sgpr_size_per_wf; // @[cta_scheduler.scala 128:51]
  assign inflight_wg_buffer_i_io_dis_controller_wg_alloc_valid = dis_controller_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 209:35 34:45]
  assign inflight_wg_buffer_i_io_dis_controller_start_alloc = dis_controller_i_io_dis_controller_start_alloc; // @[cta_scheduler.scala 207:32 35:42]
  assign inflight_wg_buffer_i_io_dis_controller_wg_dealloc_valid = dis_controller_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 210:37 36:47]
  assign inflight_wg_buffer_i_io_dis_controller_wg_rejected_valid = dis_controller_i_io_dis_controller_wg_rejected_valid
    ; // @[cta_scheduler.scala 211:38 37:48]
  assign inflight_wg_buffer_i_io_allocator_wg_id_out = allocator_neo_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 38:35 91:25]
  assign inflight_wg_buffer_i_io_gpu_interface_dealloc_wg_id = gpu_interface_i_io_gpu_interface_dealloc_wg_id; // @[cta_scheduler.scala 166:33 39:43]
  assign gpu_interface_i_clock = clock;
  assign gpu_interface_i_reset = reset;
  assign gpu_interface_i_io_inflight_wg_buffer_gpu_valid = inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_valid; // @[cta_scheduler.scala 145:34 47:44]
  assign gpu_interface_i_io_inflight_wg_buffer_gpu_wf_size = inflight_wg_buffer_i_io_inflight_wg_buffer_gpu_wf_size; // @[cta_scheduler.scala 148:36 50:46]
  assign gpu_interface_i_io_inflight_wg_buffer_start_pc = inflight_wg_buffer_i_io_inflight_wg_buffer_start_pc; // @[cta_scheduler.scala 149:33 51:43]
  assign gpu_interface_i_io_inflight_wg_buffer_gpu_vgpr_size_per_wf = inflight_wg_buffer_gpu_vgpr_size_per_wf[11:0]; // @[cta_scheduler.scala 153:64]
  assign gpu_interface_i_io_inflight_wg_buffer_gpu_sgpr_size_per_wf = inflight_wg_buffer_gpu_sgpr_size_per_wf[11:0]; // @[cta_scheduler.scala 154:64]
  assign gpu_interface_i_io_allocator_wg_id_out = allocator_neo_i_io_allocator_wg_id_out; // @[cta_scheduler.scala 38:35 91:25]
  assign gpu_interface_i_io_allocator_cu_id_out = allocator_neo_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 52:35 92:25]
  assign gpu_interface_i_io_allocator_wf_count = allocator_neo_i_io_allocator_wf_count; // @[cta_scheduler.scala 53:34 93:24]
  assign gpu_interface_i_io_allocator_vgpr_start_out = allocator_neo_i_io_allocator_vgpr_start_out; // @[cta_scheduler.scala 54:40 97:30]
  assign gpu_interface_i_io_allocator_sgpr_start_out = allocator_neo_i_io_allocator_sgpr_start_out; // @[cta_scheduler.scala 55:40 98:30]
  assign gpu_interface_i_io_allocator_lds_start_out = allocator_neo_i_io_allocator_lds_start_out; // @[cta_scheduler.scala 56:39 99:29]
  assign gpu_interface_i_io_dis_controller_wg_alloc_valid = dis_controller_i_io_dis_controller_wg_alloc_valid; // @[cta_scheduler.scala 209:35 34:45]
  assign gpu_interface_i_io_dis_controller_wg_dealloc_valid = dis_controller_i_io_dis_controller_wg_dealloc_valid; // @[cta_scheduler.scala 210:37 36:47]
  assign gpu_interface_i_io_cu2dispatch_wf_done = io_cu2dispatch_wf_done; // @[cta_scheduler.scala 175:44]
  assign gpu_interface_i_io_cu2dispatch_wf_tag_done_0 = io_cu2dispatch_wf_tag_done_0; // @[cta_scheduler.scala 176:48]
  assign gpu_interface_i_io_cu2dispatch_wf_tag_done_1 = io_cu2dispatch_wf_tag_done_1; // @[cta_scheduler.scala 176:48]
  assign gpu_interface_i_io_cu2dispatch_ready_for_dispatch_0 = io_cu2dispatch_ready_for_dispatch_0; // @[cta_scheduler.scala 177:55]
  assign gpu_interface_i_io_cu2dispatch_ready_for_dispatch_1 = io_cu2dispatch_ready_for_dispatch_1; // @[cta_scheduler.scala 177:55]
  assign dis_controller_i_clock = clock;
  assign dis_controller_i_reset = reset;
  assign dis_controller_i_io_inflight_wg_buffer_alloc_valid = inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_valid; // @[cta_scheduler.scala 138:36 40:46]
  assign dis_controller_i_io_inflight_wg_buffer_alloc_available =
    inflight_wg_buffer_i_io_inflight_wg_buffer_alloc_available; // @[cta_scheduler.scala 139:40 41:50]
  assign dis_controller_i_io_allocator_cu_valid = allocator_neo_i_io_allocator_cu_valid; // @[cta_scheduler.scala 81:34 89:24]
  assign dis_controller_i_io_allocator_cu_rejected = allocator_neo_i_io_allocator_cu_rejected; // @[cta_scheduler.scala 82:37 90:27]
  assign dis_controller_i_io_allocator_cu_id_out = allocator_neo_i_io_allocator_cu_id_out; // @[cta_scheduler.scala 52:35 92:25]
  assign dis_controller_i_io_grt_wg_alloc_done = top_resource_table_i_io_grt_wg_alloc_done; // @[cta_scheduler.scala 188:23 70:33]
  assign dis_controller_i_io_grt_wg_dealloc_done = top_resource_table_i_io_grt_wg_dealloc_done; // @[cta_scheduler.scala 191:25 73:35]
  assign dis_controller_i_io_grt_wg_alloc_cu_id = top_resource_table_i_io_grt_wg_alloc_cu_id; // @[cta_scheduler.scala 190:24 72:34]
  assign dis_controller_i_io_grt_wg_dealloc_cu_id = top_resource_table_i_io_grt_wg_dealloc_cu_id; // @[cta_scheduler.scala 193:26 75:36]
  assign dis_controller_i_io_gpu_interface_alloc_available = gpu_interface_i_io_gpu_interface_alloc_available; // @[cta_scheduler.scala 163:35 57:45]
  assign dis_controller_i_io_gpu_interface_dealloc_available = gpu_interface_i_io_gpu_interface_dealloc_available; // @[cta_scheduler.scala 164:37 58:47]
  assign dis_controller_i_io_gpu_interface_cu_id = gpu_interface_i_io_gpu_interface_cu_id; // @[cta_scheduler.scala 165:25 59:35]
endmodule
module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [4:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [4:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] ram [0:7]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[4:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module wf_done_interface_single(
  input        clock,
  input        reset,
  input        io_wf_done,
  input  [4:0] io_wf_done_wg_id,
  input        io_host_wf_done_ready,
  output       io_host_wf_done_valid,
  output [4:0] io_host_wf_done_wg_id
);
  wire  buffer_clock; // @[wf_done_interface.scala 51:24]
  wire  buffer_reset; // @[wf_done_interface.scala 51:24]
  wire  buffer_io_enq_ready; // @[wf_done_interface.scala 51:24]
  wire  buffer_io_enq_valid; // @[wf_done_interface.scala 51:24]
  wire [4:0] buffer_io_enq_bits; // @[wf_done_interface.scala 51:24]
  wire  buffer_io_deq_ready; // @[wf_done_interface.scala 51:24]
  wire  buffer_io_deq_valid; // @[wf_done_interface.scala 51:24]
  wire [4:0] buffer_io_deq_bits; // @[wf_done_interface.scala 51:24]
  Queue buffer ( // @[wf_done_interface.scala 51:24]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .io_enq_ready(buffer_io_enq_ready),
    .io_enq_valid(buffer_io_enq_valid),
    .io_enq_bits(buffer_io_enq_bits),
    .io_deq_ready(buffer_io_deq_ready),
    .io_deq_valid(buffer_io_deq_valid),
    .io_deq_bits(buffer_io_deq_bits)
  );
  assign io_host_wf_done_valid = buffer_io_deq_valid; // @[wf_done_interface.scala 55:26]
  assign io_host_wf_done_wg_id = buffer_io_deq_bits; // @[wf_done_interface.scala 54:26]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_io_enq_valid = io_wf_done; // @[wf_done_interface.scala 53:24]
  assign buffer_io_enq_bits = io_wf_done_wg_id; // @[wf_done_interface.scala 52:23]
  assign buffer_io_deq_ready = io_host_wf_done_ready; // @[wf_done_interface.scala 56:24]
endmodule
module CTAinterface(
  input         clock,
  input         reset,
  output        io_host2CTA_ready,
  input         io_host2CTA_valid,
  input  [4:0]  io_host2CTA_bits_host_wg_id,
  input  [2:0]  io_host2CTA_bits_host_num_wf,
  input  [9:0]  io_host2CTA_bits_host_wf_size,
  input  [31:0] io_host2CTA_bits_host_start_pc,
  input  [12:0] io_host2CTA_bits_host_vgpr_size_total,
  input  [12:0] io_host2CTA_bits_host_sgpr_size_total,
  input  [12:0] io_host2CTA_bits_host_lds_size_total,
  input  [10:0] io_host2CTA_bits_host_gds_size_total,
  input  [12:0] io_host2CTA_bits_host_vgpr_size_per_wf,
  input  [12:0] io_host2CTA_bits_host_sgpr_size_per_wf,
  input         io_CTA2host_ready,
  output        io_CTA2host_valid,
  output [4:0]  io_CTA2host_bits_inflight_wg_buffer_host_wf_done_wg_id,
  input         io_CTA2warp_0_ready,
  output        io_CTA2warp_0_valid,
  output [2:0]  io_CTA2warp_0_bits_dispatch2cu_wg_wf_count,
  output [9:0]  io_CTA2warp_0_bits_dispatch2cu_wf_size_dispatch,
  output [12:0] io_CTA2warp_0_bits_dispatch2cu_sgpr_base_dispatch,
  output [12:0] io_CTA2warp_0_bits_dispatch2cu_vgpr_base_dispatch,
  output [4:0]  io_CTA2warp_0_bits_dispatch2cu_wf_tag_dispatch,
  output [12:0] io_CTA2warp_0_bits_dispatch2cu_lds_base_dispatch,
  output [31:0] io_CTA2warp_0_bits_dispatch2cu_start_pc_dispatch,
  input         io_CTA2warp_1_ready,
  output        io_CTA2warp_1_valid,
  output [2:0]  io_CTA2warp_1_bits_dispatch2cu_wg_wf_count,
  output [9:0]  io_CTA2warp_1_bits_dispatch2cu_wf_size_dispatch,
  output [12:0] io_CTA2warp_1_bits_dispatch2cu_sgpr_base_dispatch,
  output [12:0] io_CTA2warp_1_bits_dispatch2cu_vgpr_base_dispatch,
  output [4:0]  io_CTA2warp_1_bits_dispatch2cu_wf_tag_dispatch,
  output [12:0] io_CTA2warp_1_bits_dispatch2cu_lds_base_dispatch,
  output [31:0] io_CTA2warp_1_bits_dispatch2cu_start_pc_dispatch,
  input         io_warp2CTA_0_valid,
  input  [4:0]  io_warp2CTA_0_bits_cu2dispatch_wf_tag_done,
  input         io_warp2CTA_1_valid,
  input  [4:0]  io_warp2CTA_1_bits_cu2dispatch_wf_tag_done
);
  wire  cta_sche_clock; // @[GPGPU_top.scala 46:22]
  wire  cta_sche_reset; // @[GPGPU_top.scala 46:22]
  wire  cta_sche_io_host_wg_valid; // @[GPGPU_top.scala 46:22]
  wire [4:0] cta_sche_io_host_wg_id; // @[GPGPU_top.scala 46:22]
  wire [2:0] cta_sche_io_host_num_wf; // @[GPGPU_top.scala 46:22]
  wire [9:0] cta_sche_io_host_wf_size; // @[GPGPU_top.scala 46:22]
  wire [31:0] cta_sche_io_host_start_pc; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_host_vgpr_size_total; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_host_sgpr_size_total; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_host_lds_size_total; // @[GPGPU_top.scala 46:22]
  wire [10:0] cta_sche_io_host_gds_size_total; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_host_vgpr_size_per_wf; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_host_sgpr_size_per_wf; // @[GPGPU_top.scala 46:22]
  wire  cta_sche_io_inflight_wg_buffer_host_rcvd_ack; // @[GPGPU_top.scala 46:22]
  wire  cta_sche_io_inflight_wg_buffer_host_wf_done; // @[GPGPU_top.scala 46:22]
  wire [4:0] cta_sche_io_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 46:22]
  wire [1:0] cta_sche_io_dispatch2cu_wf_dispatch; // @[GPGPU_top.scala 46:22]
  wire [2:0] cta_sche_io_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 46:22]
  wire [9:0] cta_sche_io_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 46:22]
  wire [4:0] cta_sche_io_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 46:22]
  wire [12:0] cta_sche_io_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 46:22]
  wire [31:0] cta_sche_io_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 46:22]
  wire [1:0] cta_sche_io_cu2dispatch_wf_done; // @[GPGPU_top.scala 46:22]
  wire [4:0] cta_sche_io_cu2dispatch_wf_tag_done_0; // @[GPGPU_top.scala 46:22]
  wire [4:0] cta_sche_io_cu2dispatch_wf_tag_done_1; // @[GPGPU_top.scala 46:22]
  wire  cta_sche_io_cu2dispatch_ready_for_dispatch_0; // @[GPGPU_top.scala 46:22]
  wire  cta_sche_io_cu2dispatch_ready_for_dispatch_1; // @[GPGPU_top.scala 46:22]
  wire  wf_done_interface_clock; // @[GPGPU_top.scala 60:31]
  wire  wf_done_interface_reset; // @[GPGPU_top.scala 60:31]
  wire  wf_done_interface_io_wf_done; // @[GPGPU_top.scala 60:31]
  wire [4:0] wf_done_interface_io_wf_done_wg_id; // @[GPGPU_top.scala 60:31]
  wire  wf_done_interface_io_host_wf_done_ready; // @[GPGPU_top.scala 60:31]
  wire  wf_done_interface_io_host_wf_done_valid; // @[GPGPU_top.scala 60:31]
  wire [4:0] wf_done_interface_io_host_wf_done_wg_id; // @[GPGPU_top.scala 60:31]
  cta_scheduler cta_sche ( // @[GPGPU_top.scala 46:22]
    .clock(cta_sche_clock),
    .reset(cta_sche_reset),
    .io_host_wg_valid(cta_sche_io_host_wg_valid),
    .io_host_wg_id(cta_sche_io_host_wg_id),
    .io_host_num_wf(cta_sche_io_host_num_wf),
    .io_host_wf_size(cta_sche_io_host_wf_size),
    .io_host_start_pc(cta_sche_io_host_start_pc),
    .io_host_vgpr_size_total(cta_sche_io_host_vgpr_size_total),
    .io_host_sgpr_size_total(cta_sche_io_host_sgpr_size_total),
    .io_host_lds_size_total(cta_sche_io_host_lds_size_total),
    .io_host_gds_size_total(cta_sche_io_host_gds_size_total),
    .io_host_vgpr_size_per_wf(cta_sche_io_host_vgpr_size_per_wf),
    .io_host_sgpr_size_per_wf(cta_sche_io_host_sgpr_size_per_wf),
    .io_inflight_wg_buffer_host_rcvd_ack(cta_sche_io_inflight_wg_buffer_host_rcvd_ack),
    .io_inflight_wg_buffer_host_wf_done(cta_sche_io_inflight_wg_buffer_host_wf_done),
    .io_inflight_wg_buffer_host_wf_done_wg_id(cta_sche_io_inflight_wg_buffer_host_wf_done_wg_id),
    .io_dispatch2cu_wf_dispatch(cta_sche_io_dispatch2cu_wf_dispatch),
    .io_dispatch2cu_wg_wf_count(cta_sche_io_dispatch2cu_wg_wf_count),
    .io_dispatch2cu_wf_size_dispatch(cta_sche_io_dispatch2cu_wf_size_dispatch),
    .io_dispatch2cu_sgpr_base_dispatch(cta_sche_io_dispatch2cu_sgpr_base_dispatch),
    .io_dispatch2cu_vgpr_base_dispatch(cta_sche_io_dispatch2cu_vgpr_base_dispatch),
    .io_dispatch2cu_wf_tag_dispatch(cta_sche_io_dispatch2cu_wf_tag_dispatch),
    .io_dispatch2cu_lds_base_dispatch(cta_sche_io_dispatch2cu_lds_base_dispatch),
    .io_dispatch2cu_start_pc_dispatch(cta_sche_io_dispatch2cu_start_pc_dispatch),
    .io_cu2dispatch_wf_done(cta_sche_io_cu2dispatch_wf_done),
    .io_cu2dispatch_wf_tag_done_0(cta_sche_io_cu2dispatch_wf_tag_done_0),
    .io_cu2dispatch_wf_tag_done_1(cta_sche_io_cu2dispatch_wf_tag_done_1),
    .io_cu2dispatch_ready_for_dispatch_0(cta_sche_io_cu2dispatch_ready_for_dispatch_0),
    .io_cu2dispatch_ready_for_dispatch_1(cta_sche_io_cu2dispatch_ready_for_dispatch_1)
  );
  wf_done_interface_single wf_done_interface ( // @[GPGPU_top.scala 60:31]
    .clock(wf_done_interface_clock),
    .reset(wf_done_interface_reset),
    .io_wf_done(wf_done_interface_io_wf_done),
    .io_wf_done_wg_id(wf_done_interface_io_wf_done_wg_id),
    .io_host_wf_done_ready(wf_done_interface_io_host_wf_done_ready),
    .io_host_wf_done_valid(wf_done_interface_io_host_wf_done_valid),
    .io_host_wf_done_wg_id(wf_done_interface_io_host_wf_done_wg_id)
  );
  assign io_host2CTA_ready = cta_sche_io_inflight_wg_buffer_host_rcvd_ack; // @[GPGPU_top.scala 58:20]
  assign io_CTA2host_valid = wf_done_interface_io_host_wf_done_valid; // @[GPGPU_top.scala 65:20]
  assign io_CTA2host_bits_inflight_wg_buffer_host_wf_done_wg_id = wf_done_interface_io_host_wf_done_wg_id; // @[GPGPU_top.scala 64:57]
  assign io_CTA2warp_0_valid = cta_sche_io_dispatch2cu_wf_dispatch[0]; // @[GPGPU_top.scala 70:62]
  assign io_CTA2warp_0_bits_dispatch2cu_wg_wf_count = cta_sche_io_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 71:48]
  assign io_CTA2warp_0_bits_dispatch2cu_wf_size_dispatch = cta_sche_io_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 72:56]
  assign io_CTA2warp_0_bits_dispatch2cu_sgpr_base_dispatch = cta_sche_io_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 73:56]
  assign io_CTA2warp_0_bits_dispatch2cu_vgpr_base_dispatch = cta_sche_io_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 74:56]
  assign io_CTA2warp_0_bits_dispatch2cu_wf_tag_dispatch = cta_sche_io_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 75:56]
  assign io_CTA2warp_0_bits_dispatch2cu_lds_base_dispatch = cta_sche_io_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 76:56]
  assign io_CTA2warp_0_bits_dispatch2cu_start_pc_dispatch = cta_sche_io_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 77:56]
  assign io_CTA2warp_1_valid = cta_sche_io_dispatch2cu_wf_dispatch[1]; // @[GPGPU_top.scala 70:62]
  assign io_CTA2warp_1_bits_dispatch2cu_wg_wf_count = cta_sche_io_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 71:48]
  assign io_CTA2warp_1_bits_dispatch2cu_wf_size_dispatch = cta_sche_io_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 72:56]
  assign io_CTA2warp_1_bits_dispatch2cu_sgpr_base_dispatch = cta_sche_io_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 73:56]
  assign io_CTA2warp_1_bits_dispatch2cu_vgpr_base_dispatch = cta_sche_io_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 74:56]
  assign io_CTA2warp_1_bits_dispatch2cu_wf_tag_dispatch = cta_sche_io_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 75:56]
  assign io_CTA2warp_1_bits_dispatch2cu_lds_base_dispatch = cta_sche_io_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 76:56]
  assign io_CTA2warp_1_bits_dispatch2cu_start_pc_dispatch = cta_sche_io_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 77:56]
  assign cta_sche_clock = clock;
  assign cta_sche_reset = reset;
  assign cta_sche_io_host_wg_valid = io_host2CTA_valid; // @[GPGPU_top.scala 47:37]
  assign cta_sche_io_host_wg_id = io_host2CTA_bits_host_wg_id; // @[GPGPU_top.scala 48:37]
  assign cta_sche_io_host_num_wf = io_host2CTA_bits_host_num_wf; // @[GPGPU_top.scala 49:37]
  assign cta_sche_io_host_wf_size = io_host2CTA_bits_host_wf_size; // @[GPGPU_top.scala 50:37]
  assign cta_sche_io_host_start_pc = io_host2CTA_bits_host_start_pc; // @[GPGPU_top.scala 51:37]
  assign cta_sche_io_host_vgpr_size_total = io_host2CTA_bits_host_vgpr_size_total; // @[GPGPU_top.scala 52:37]
  assign cta_sche_io_host_sgpr_size_total = io_host2CTA_bits_host_sgpr_size_total; // @[GPGPU_top.scala 53:37]
  assign cta_sche_io_host_lds_size_total = io_host2CTA_bits_host_lds_size_total; // @[GPGPU_top.scala 54:37]
  assign cta_sche_io_host_gds_size_total = io_host2CTA_bits_host_gds_size_total; // @[GPGPU_top.scala 55:37]
  assign cta_sche_io_host_vgpr_size_per_wf = io_host2CTA_bits_host_vgpr_size_per_wf; // @[GPGPU_top.scala 56:37]
  assign cta_sche_io_host_sgpr_size_per_wf = io_host2CTA_bits_host_sgpr_size_per_wf; // @[GPGPU_top.scala 57:37]
  assign cta_sche_io_cu2dispatch_wf_done = {io_warp2CTA_1_valid,io_warp2CTA_0_valid}; // @[GPGPU_top.scala 84:56]
  assign cta_sche_io_cu2dispatch_wf_tag_done_0 = io_warp2CTA_0_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 80:43]
  assign cta_sche_io_cu2dispatch_wf_tag_done_1 = io_warp2CTA_1_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 80:43]
  assign cta_sche_io_cu2dispatch_ready_for_dispatch_0 = io_CTA2warp_0_ready; // @[GPGPU_top.scala 78:50]
  assign cta_sche_io_cu2dispatch_ready_for_dispatch_1 = io_CTA2warp_1_ready; // @[GPGPU_top.scala 78:50]
  assign wf_done_interface_clock = clock;
  assign wf_done_interface_reset = reset;
  assign wf_done_interface_io_wf_done = cta_sche_io_inflight_wg_buffer_host_wf_done; // @[GPGPU_top.scala 61:31]
  assign wf_done_interface_io_wf_done_wg_id = cta_sche_io_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 62:37]
  assign wf_done_interface_io_host_wf_done_ready = io_CTA2host_ready; // @[GPGPU_top.scala 66:42]
endmodule
module CTA2warp(
  input         clock,
  input         reset,
  output        io_CTAreq_ready,
  input         io_CTAreq_valid,
  input  [2:0]  io_CTAreq_bits_dispatch2cu_wg_wf_count,
  input  [9:0]  io_CTAreq_bits_dispatch2cu_wf_size_dispatch,
  input  [12:0] io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch,
  input  [12:0] io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch,
  input  [4:0]  io_CTAreq_bits_dispatch2cu_wf_tag_dispatch,
  input  [12:0] io_CTAreq_bits_dispatch2cu_lds_base_dispatch,
  input  [31:0] io_CTAreq_bits_dispatch2cu_start_pc_dispatch,
  output        io_CTArsp_valid,
  output [4:0]  io_CTArsp_bits_cu2dispatch_wf_tag_done,
  output        io_warpReq_valid,
  output [2:0]  io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count,
  output [9:0]  io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch,
  output [12:0] io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch,
  output [12:0] io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch,
  output [4:0]  io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch,
  output [12:0] io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch,
  output [31:0] io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch,
  output [1:0]  io_warpReq_bits_wid,
  output        io_warpRsp_ready,
  input         io_warpRsp_valid,
  input  [1:0]  io_warpRsp_bits_wid,
  input  [1:0]  io_wg_id_lookup,
  output [4:0]  io_wg_id_tag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] idx_using; // @[CTA2warp.scala 36:26]
  reg [4:0] data_0; // @[CTA2warp.scala 39:17]
  reg [4:0] data_1; // @[CTA2warp.scala 39:17]
  reg [4:0] data_2; // @[CTA2warp.scala 39:17]
  reg [4:0] data_3; // @[CTA2warp.scala 39:17]
  wire [4:0] _GEN_1 = 2'h1 == io_wg_id_lookup ? data_1 : data_0; // @[CTA2warp.scala 40:{15,15}]
  wire [4:0] _GEN_2 = 2'h2 == io_wg_id_lookup ? data_2 : _GEN_1; // @[CTA2warp.scala 40:{15,15}]
  wire [3:0] _idx_next_allocate_T = ~idx_using; // @[CTA2warp.scala 41:43]
  wire [1:0] _idx_next_allocate_T_5 = _idx_next_allocate_T[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _idx_next_allocate_T_6 = _idx_next_allocate_T[1] ? 2'h1 : _idx_next_allocate_T_5; // @[Mux.scala 47:70]
  wire [1:0] idx_next_allocate = _idx_next_allocate_T[0] ? 2'h0 : _idx_next_allocate_T_6; // @[Mux.scala 47:70]
  wire [3:0] _idx_using_T = 4'h1 << idx_next_allocate; // @[CTA2warp.scala 45:32]
  wire  _idx_using_T_1 = io_CTAreq_ready & io_CTAreq_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _idx_using_T_3 = _idx_using_T_1 ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _idx_using_T_4 = _idx_using_T & _idx_using_T_3; // @[CTA2warp.scala 45:60]
  wire [3:0] _idx_using_T_5 = idx_using | _idx_using_T_4; // @[CTA2warp.scala 45:25]
  wire  _idx_using_T_6 = io_warpRsp_ready & io_warpRsp_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _idx_using_T_8 = _idx_using_T_6 ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _idx_using_T_9 = 4'h1 << io_warpRsp_bits_wid; // @[CTA2warp.scala 45:148]
  wire [3:0] _idx_using_T_10 = _idx_using_T_8 & _idx_using_T_9; // @[CTA2warp.scala 45:141]
  wire [3:0] _idx_using_T_11 = ~_idx_using_T_10; // @[CTA2warp.scala 45:97]
  wire [3:0] _idx_using_T_12 = _idx_using_T_5 & _idx_using_T_11; // @[CTA2warp.scala 45:94]
  wire [4:0] _GEN_13 = 2'h1 == io_warpRsp_bits_wid ? data_1 : data_0; // @[CTA2warp.scala 53:{41,41}]
  wire [4:0] _GEN_14 = 2'h2 == io_warpRsp_bits_wid ? data_2 : _GEN_13; // @[CTA2warp.scala 53:{41,41}]
  assign io_CTAreq_ready = ~(&idx_using); // @[CTA2warp.scala 38:21]
  assign io_CTArsp_valid = io_warpRsp_valid; // @[CTA2warp.scala 54:18]
  assign io_CTArsp_bits_cu2dispatch_wf_tag_done = 2'h3 == io_warpRsp_bits_wid ? data_3 : _GEN_14; // @[CTA2warp.scala 53:{41,41}]
  assign io_warpReq_valid = io_CTAreq_ready & io_CTAreq_valid; // @[Decoupled.scala 50:35]
  assign io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count = io_CTAreq_bits_dispatch2cu_wg_wf_count; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch = io_CTAreq_bits_dispatch2cu_wf_size_dispatch; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch = io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch = io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch = io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch = io_CTAreq_bits_dispatch2cu_lds_base_dispatch; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch = io_CTAreq_bits_dispatch2cu_start_pc_dispatch; // @[CTA2warp.scala 50:26]
  assign io_warpReq_bits_wid = _idx_next_allocate_T[0] ? 2'h0 : _idx_next_allocate_T_6; // @[Mux.scala 47:70]
  assign io_warpRsp_ready = 1'h1; // @[CTA2warp.scala 52:19]
  assign io_wg_id_tag = 2'h3 == io_wg_id_lookup ? data_3 : _GEN_2; // @[CTA2warp.scala 40:{15,15}]
  always @(posedge clock) begin
    if (reset) begin // @[CTA2warp.scala 36:26]
      idx_using <= 4'h0; // @[CTA2warp.scala 36:26]
    end else begin
      idx_using <= _idx_using_T_12; // @[CTA2warp.scala 45:12]
    end
    if (_idx_using_T_1) begin // @[CTA2warp.scala 46:24]
      if (2'h0 == idx_next_allocate) begin // @[CTA2warp.scala 47:28]
        data_0 <= io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[CTA2warp.scala 47:28]
      end
    end
    if (_idx_using_T_1) begin // @[CTA2warp.scala 46:24]
      if (2'h1 == idx_next_allocate) begin // @[CTA2warp.scala 47:28]
        data_1 <= io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[CTA2warp.scala 47:28]
      end
    end
    if (_idx_using_T_1) begin // @[CTA2warp.scala 46:24]
      if (2'h2 == idx_next_allocate) begin // @[CTA2warp.scala 47:28]
        data_2 <= io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[CTA2warp.scala 47:28]
      end
    end
    if (_idx_using_T_1) begin // @[CTA2warp.scala 46:24]
      if (2'h3 == idx_next_allocate) begin // @[CTA2warp.scala 47:28]
        data_3 <= io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[CTA2warp.scala 47:28]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idx_using = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  data_0 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  data_1 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  data_2 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  data_3 = _RAND_4[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PCcontrol(
  input         clock,
  input         reset,
  input  [31:0] io_New_PC,
  input         io_PC_replay,
  input  [1:0]  io_PC_src,
  output [31:0] io_PC_next
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pout; // @[PCcontrol.scala 13:19]
  wire [31:0] _pout_T_1 = pout + 32'h4; // @[PCcontrol.scala 19:15]
  wire [31:0] _pout_T_3 = pout - 32'h8; // @[PCcontrol.scala 23:15]
  wire [31:0] _GEN_0 = io_PC_src == 2'h3 ? _pout_T_3 : pout; // @[PCcontrol.scala 22:30 23:9 25:9]
  assign io_PC_next = pout; // @[PCcontrol.scala 27:13]
  always @(posedge clock) begin
    if (reset) begin // @[PCcontrol.scala 13:19]
      pout <= 32'h0; // @[PCcontrol.scala 13:19]
    end else if (!(io_PC_replay)) begin // @[PCcontrol.scala 16:21]
      if (io_PC_src == 2'h2) begin // @[PCcontrol.scala 18:30]
        pout <= _pout_T_1; // @[PCcontrol.scala 19:9]
      end else if (io_PC_src == 2'h1) begin // @[PCcontrol.scala 20:30]
        pout <= io_New_PC; // @[PCcontrol.scala 21:9]
      end else begin
        pout <= _GEN_0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pout = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module warp_scheduler(
  input         clock,
  input         reset,
  input         io_pc_reset,
  output        io_warpReq_ready,
  input         io_warpReq_valid,
  input  [2:0]  io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count,
  input  [9:0]  io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch,
  input  [12:0] io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch,
  input  [12:0] io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch,
  input  [4:0]  io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch,
  input  [12:0] io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch,
  input  [31:0] io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch,
  input  [1:0]  io_warpReq_bits_wid,
  output        io_warpRsp_valid,
  output [1:0]  io_warpRsp_bits_wid,
  output [1:0]  io_wg_id_lookup,
  input  [4:0]  io_wg_id_tag,
  output        io_pc_req_valid,
  output [31:0] io_pc_req_bits_addr,
  output [1:0]  io_pc_req_bits_warpid,
  input         io_pc_rsp_valid,
  input  [31:0] io_pc_rsp_bits_addr,
  input  [1:0]  io_pc_rsp_bits_warpid,
  input  [1:0]  io_pc_rsp_bits_status,
  output        io_branch_ready,
  input         io_branch_valid,
  input  [1:0]  io_branch_bits_wid,
  input         io_branch_bits_jump,
  input  [31:0] io_branch_bits_new_pc,
  output        io_warp_control_ready,
  input         io_warp_control_valid,
  input  [1:0]  io_warp_control_bits_ctrl_wid,
  input         io_warp_control_bits_ctrl_simt_stack_op,
  input         io_warp_control_bits_ctrl_barrier,
  input  [3:0]  io_scoreboard_busy,
  input  [3:0]  io_exe_busy,
  input         io_pc_ibuffer_ready_0,
  input         io_pc_ibuffer_ready_1,
  input         io_pc_ibuffer_ready_2,
  input         io_pc_ibuffer_ready_3,
  output [3:0]  io_warp_ready,
  output        io_flush_valid,
  output [1:0]  io_flush_bits,
  output        io_flushCache_valid,
  output [1:0]  io_flushCache_bits,
  output        io_CTA2csr_valid,
  output [2:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count,
  output [9:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch,
  output [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch,
  output [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch,
  output [4:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch,
  output [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch,
  output [1:0]  io_CTA2csr_bits_wid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  PCcontrol_clock; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_reset; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_io_New_PC; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_io_PC_replay; // @[warp_schedule.scala 50:50]
  wire [1:0] PCcontrol_io_PC_src; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_io_PC_next; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_1_clock; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_1_reset; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_1_io_New_PC; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_1_io_PC_replay; // @[warp_schedule.scala 50:50]
  wire [1:0] PCcontrol_1_io_PC_src; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_1_io_PC_next; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_2_clock; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_2_reset; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_2_io_New_PC; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_2_io_PC_replay; // @[warp_schedule.scala 50:50]
  wire [1:0] PCcontrol_2_io_PC_src; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_2_io_PC_next; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_3_clock; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_3_reset; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_3_io_New_PC; // @[warp_schedule.scala 50:50]
  wire  PCcontrol_3_io_PC_replay; // @[warp_schedule.scala 50:50]
  wire [1:0] PCcontrol_3_io_PC_src; // @[warp_schedule.scala 50:50]
  wire [31:0] PCcontrol_3_io_PC_next; // @[warp_schedule.scala 50:50]
  wire  _warp_end_T = io_warp_control_ready & io_warp_control_valid; // @[Decoupled.scala 50:35]
  wire  warp_end = _warp_end_T & io_warp_control_bits_ctrl_simt_stack_op; // @[warp_schedule.scala 31:38]
  wire  _io_branch_ready_T = ~io_flushCache_valid; // @[warp_schedule.scala 34:21]
  wire  _io_warp_control_ready_T = io_branch_ready & io_branch_valid; // @[Decoupled.scala 50:35]
  wire  _io_flush_valid_T_1 = _io_warp_control_ready_T & io_branch_bits_jump; // @[warp_schedule.scala 45:36]
  wire  _io_flushCache_valid_T_1 = io_pc_rsp_valid & io_pc_rsp_bits_status[0]; // @[warp_schedule.scala 47:39]
  reg [1:0] current_warp; // @[warp_schedule.scala 65:27]
  reg [3:0] warp_active; // @[warp_schedule.scala 113:26]
  wire  pc_ready_0 = io_pc_ibuffer_ready_0 & warp_active[0]; // @[warp_schedule.scala 122:42]
  wire  pc_ready_1 = io_pc_ibuffer_ready_1 & warp_active[1]; // @[warp_schedule.scala 122:42]
  wire  pc_ready_2 = io_pc_ibuffer_ready_2 & warp_active[2]; // @[warp_schedule.scala 122:42]
  wire  pc_ready_3 = io_pc_ibuffer_ready_3 & warp_active[3]; // @[warp_schedule.scala 122:42]
  wire [1:0] _GEN_102 = pc_ready_3 ? 2'h3 : current_warp; // @[warp_schedule.scala 124:{22,32}]
  wire [1:0] _GEN_103 = pc_ready_2 ? 2'h2 : _GEN_102; // @[warp_schedule.scala 124:{22,32}]
  wire [1:0] _GEN_104 = pc_ready_1 ? 2'h1 : _GEN_103; // @[warp_schedule.scala 124:{22,32}]
  wire [1:0] next_warp = pc_ready_0 ? 2'h0 : _GEN_104; // @[warp_schedule.scala 124:{22,32}]
  wire  _GEN_1 = 2'h1 == next_warp ? pc_ready_1 : pc_ready_0; // @[warp_schedule.scala 68:{56,56}]
  wire  _GEN_2 = 2'h2 == next_warp ? pc_ready_2 : _GEN_1; // @[warp_schedule.scala 68:{56,56}]
  wire  _GEN_3 = 2'h3 == next_warp ? pc_ready_3 : _GEN_2; // @[warp_schedule.scala 68:{56,56}]
  wire  _GEN_4 = 2'h0 == next_warp ? ~_GEN_3 : 1'h1; // @[warp_schedule.scala 59:18 68:{33,33}]
  wire  _GEN_5 = 2'h1 == next_warp ? ~_GEN_3 : 1'h1; // @[warp_schedule.scala 59:18 68:{33,33}]
  wire  _GEN_6 = 2'h2 == next_warp ? ~_GEN_3 : 1'h1; // @[warp_schedule.scala 59:18 68:{33,33}]
  wire  _GEN_7 = 2'h3 == next_warp ? ~_GEN_3 : 1'h1; // @[warp_schedule.scala 59:18 68:{33,33}]
  wire [1:0] _GEN_8 = 2'h0 == next_warp ? 2'h2 : 2'h0; // @[warp_schedule.scala 60:15 69:{30,30}]
  wire [1:0] _GEN_9 = 2'h1 == next_warp ? 2'h2 : 2'h0; // @[warp_schedule.scala 60:15 69:{30,30}]
  wire [1:0] _GEN_10 = 2'h2 == next_warp ? 2'h2 : 2'h0; // @[warp_schedule.scala 60:15 69:{30,30}]
  wire [1:0] _GEN_11 = 2'h3 == next_warp ? 2'h2 : 2'h0; // @[warp_schedule.scala 60:15 69:{30,30}]
  wire [31:0] pcControl_0_PC_next = PCcontrol_io_PC_next; // @[warp_schedule.scala 50:{24,24}]
  wire [31:0] pcControl_1_PC_next = PCcontrol_1_io_PC_next; // @[warp_schedule.scala 50:{24,24}]
  wire [31:0] _GEN_13 = 2'h1 == next_warp ? pcControl_1_PC_next : pcControl_0_PC_next; // @[warp_schedule.scala 72:{22,22}]
  wire [31:0] pcControl_2_PC_next = PCcontrol_2_io_PC_next; // @[warp_schedule.scala 50:{24,24}]
  wire [31:0] _GEN_14 = 2'h2 == next_warp ? pcControl_2_PC_next : _GEN_13; // @[warp_schedule.scala 72:{22,22}]
  wire [31:0] pcControl_3_PC_next = PCcontrol_3_io_PC_next; // @[warp_schedule.scala 50:{24,24}]
  reg [3:0] warp_bar_cur_0; // @[warp_schedule.scala 77:27]
  reg [3:0] warp_bar_cur_1; // @[warp_schedule.scala 77:27]
  reg [3:0] warp_bar_cur_2; // @[warp_schedule.scala 77:27]
  reg [3:0] warp_bar_cur_3; // @[warp_schedule.scala 77:27]
  reg [3:0] warp_bar_exp_0; // @[warp_schedule.scala 78:27]
  reg [3:0] warp_bar_exp_1; // @[warp_schedule.scala 78:27]
  reg [3:0] warp_bar_exp_2; // @[warp_schedule.scala 78:27]
  reg [3:0] warp_bar_exp_3; // @[warp_schedule.scala 78:27]
  reg  warp_bar_lock_0; // @[warp_schedule.scala 81:28]
  reg  warp_bar_lock_1; // @[warp_schedule.scala 81:28]
  reg  warp_bar_lock_2; // @[warp_schedule.scala 81:28]
  reg  warp_bar_lock_3; // @[warp_schedule.scala 81:28]
  wire [1:0] new_wg_id = io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch[4:3]; // @[warp_schedule.scala 82:68]
  wire [1:0] end_wg_id = io_wg_id_tag[4:3]; // @[warp_schedule.scala 85:29]
  wire [2:0] end_wf_id = io_wg_id_tag[2:0]; // @[warp_schedule.scala 86:29]
  reg [3:0] warp_bar_data; // @[warp_schedule.scala 87:28]
  reg [3:0] warp_bar_belong_0; // @[warp_schedule.scala 88:30]
  reg [3:0] warp_bar_belong_1; // @[warp_schedule.scala 88:30]
  reg [3:0] warp_bar_belong_2; // @[warp_schedule.scala 88:30]
  reg [3:0] warp_bar_belong_3; // @[warp_schedule.scala 88:30]
  wire  _T_4 = io_warpReq_ready & io_warpReq_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _warp_bar_belong_T = 4'h1 << io_warpReq_bits_wid; // @[warp_schedule.scala 91:66]
  wire [3:0] _GEN_17 = 2'h1 == new_wg_id ? warp_bar_belong_1 : warp_bar_belong_0; // @[warp_schedule.scala 91:{60,60}]
  wire [3:0] _GEN_18 = 2'h2 == new_wg_id ? warp_bar_belong_2 : _GEN_17; // @[warp_schedule.scala 91:{60,60}]
  wire [3:0] _GEN_19 = 2'h3 == new_wg_id ? warp_bar_belong_3 : _GEN_18; // @[warp_schedule.scala 91:{60,60}]
  wire [3:0] _warp_bar_belong_T_1 = _GEN_19 | _warp_bar_belong_T; // @[warp_schedule.scala 91:60]
  wire [3:0] _GEN_20 = 2'h0 == new_wg_id ? _warp_bar_belong_T_1 : warp_bar_belong_0; // @[warp_schedule.scala 88:30 91:{31,31}]
  wire [3:0] _GEN_21 = 2'h1 == new_wg_id ? _warp_bar_belong_T_1 : warp_bar_belong_1; // @[warp_schedule.scala 88:30 91:{31,31}]
  wire [3:0] _GEN_22 = 2'h2 == new_wg_id ? _warp_bar_belong_T_1 : warp_bar_belong_2; // @[warp_schedule.scala 88:30 91:{31,31}]
  wire [3:0] _GEN_23 = 2'h3 == new_wg_id ? _warp_bar_belong_T_1 : warp_bar_belong_3; // @[warp_schedule.scala 88:30 91:{31,31}]
  wire  _GEN_25 = 2'h1 == new_wg_id ? warp_bar_lock_1 : warp_bar_lock_0; // @[warp_schedule.scala 92:{10,10}]
  wire  _GEN_26 = 2'h2 == new_wg_id ? warp_bar_lock_2 : _GEN_25; // @[warp_schedule.scala 92:{10,10}]
  wire  _GEN_27 = 2'h3 == new_wg_id ? warp_bar_lock_3 : _GEN_26; // @[warp_schedule.scala 92:{10,10}]
  wire [2:0] _warp_bar_exp_T_2 = 3'h4 - io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count; // @[warp_schedule.scala 93:96]
  wire [3:0] _warp_bar_exp_T_3 = 4'hf >> _warp_bar_exp_T_2; // @[warp_schedule.scala 93:67]
  wire [3:0] _GEN_28 = 2'h0 == new_wg_id ? _warp_bar_exp_T_3 : warp_bar_exp_0; // @[warp_schedule.scala 78:27 93:{30,30}]
  wire [3:0] _GEN_29 = 2'h1 == new_wg_id ? _warp_bar_exp_T_3 : warp_bar_exp_1; // @[warp_schedule.scala 78:27 93:{30,30}]
  wire [3:0] _GEN_30 = 2'h2 == new_wg_id ? _warp_bar_exp_T_3 : warp_bar_exp_2; // @[warp_schedule.scala 78:27 93:{30,30}]
  wire [3:0] _GEN_31 = 2'h3 == new_wg_id ? _warp_bar_exp_T_3 : warp_bar_exp_3; // @[warp_schedule.scala 78:27 93:{30,30}]
  wire [3:0] _GEN_32 = 2'h0 == new_wg_id ? 4'h0 : warp_bar_cur_0; // @[warp_schedule.scala 77:27 94:{30,30}]
  wire [3:0] _GEN_33 = 2'h1 == new_wg_id ? 4'h0 : warp_bar_cur_1; // @[warp_schedule.scala 77:27 94:{30,30}]
  wire [3:0] _GEN_34 = 2'h2 == new_wg_id ? 4'h0 : warp_bar_cur_2; // @[warp_schedule.scala 77:27 94:{30,30}]
  wire [3:0] _GEN_35 = 2'h3 == new_wg_id ? 4'h0 : warp_bar_cur_3; // @[warp_schedule.scala 77:27 94:{30,30}]
  wire [3:0] _GEN_36 = ~_GEN_27 ? _GEN_28 : warp_bar_exp_0; // @[warp_schedule.scala 78:27 92:36]
  wire [3:0] _GEN_37 = ~_GEN_27 ? _GEN_29 : warp_bar_exp_1; // @[warp_schedule.scala 78:27 92:36]
  wire [3:0] _GEN_38 = ~_GEN_27 ? _GEN_30 : warp_bar_exp_2; // @[warp_schedule.scala 78:27 92:36]
  wire [3:0] _GEN_39 = ~_GEN_27 ? _GEN_31 : warp_bar_exp_3; // @[warp_schedule.scala 78:27 92:36]
  wire [3:0] _GEN_40 = ~_GEN_27 ? _GEN_32 : warp_bar_cur_0; // @[warp_schedule.scala 77:27 92:36]
  wire [3:0] _GEN_41 = ~_GEN_27 ? _GEN_33 : warp_bar_cur_1; // @[warp_schedule.scala 77:27 92:36]
  wire [3:0] _GEN_42 = ~_GEN_27 ? _GEN_34 : warp_bar_cur_2; // @[warp_schedule.scala 77:27 92:36]
  wire [3:0] _GEN_43 = ~_GEN_27 ? _GEN_35 : warp_bar_cur_3; // @[warp_schedule.scala 77:27 92:36]
  wire [3:0] _GEN_44 = _T_4 ? _GEN_20 : warp_bar_belong_0; // @[warp_schedule.scala 90:24 88:30]
  wire [3:0] _GEN_45 = _T_4 ? _GEN_21 : warp_bar_belong_1; // @[warp_schedule.scala 90:24 88:30]
  wire [3:0] _GEN_46 = _T_4 ? _GEN_22 : warp_bar_belong_2; // @[warp_schedule.scala 90:24 88:30]
  wire [3:0] _GEN_47 = _T_4 ? _GEN_23 : warp_bar_belong_3; // @[warp_schedule.scala 90:24 88:30]
  wire [3:0] _GEN_48 = _T_4 ? _GEN_36 : warp_bar_exp_0; // @[warp_schedule.scala 90:24 78:27]
  wire [3:0] _GEN_49 = _T_4 ? _GEN_37 : warp_bar_exp_1; // @[warp_schedule.scala 90:24 78:27]
  wire [3:0] _GEN_50 = _T_4 ? _GEN_38 : warp_bar_exp_2; // @[warp_schedule.scala 90:24 78:27]
  wire [3:0] _GEN_51 = _T_4 ? _GEN_39 : warp_bar_exp_3; // @[warp_schedule.scala 90:24 78:27]
  wire [3:0] _GEN_52 = _T_4 ? _GEN_40 : warp_bar_cur_0; // @[warp_schedule.scala 90:24 77:27]
  wire [3:0] _GEN_53 = _T_4 ? _GEN_41 : warp_bar_cur_1; // @[warp_schedule.scala 90:24 77:27]
  wire [3:0] _GEN_54 = _T_4 ? _GEN_42 : warp_bar_cur_2; // @[warp_schedule.scala 90:24 77:27]
  wire [3:0] _GEN_55 = _T_4 ? _GEN_43 : warp_bar_cur_3; // @[warp_schedule.scala 90:24 77:27]
  wire [7:0] _warp_bar_exp_T_4 = 8'h1 << end_wf_id; // @[warp_schedule.scala 98:62]
  wire [7:0] _warp_bar_exp_T_5 = ~_warp_bar_exp_T_4; // @[warp_schedule.scala 98:57]
  wire [3:0] _GEN_57 = 2'h1 == end_wg_id ? warp_bar_exp_1 : warp_bar_exp_0; // @[warp_schedule.scala 98:{54,54}]
  wire [3:0] _GEN_58 = 2'h2 == end_wg_id ? warp_bar_exp_2 : _GEN_57; // @[warp_schedule.scala 98:{54,54}]
  wire [3:0] _GEN_59 = 2'h3 == end_wg_id ? warp_bar_exp_3 : _GEN_58; // @[warp_schedule.scala 98:{54,54}]
  wire [7:0] _GEN_197 = {{4'd0}, _GEN_59}; // @[warp_schedule.scala 98:54]
  wire [7:0] _warp_bar_exp_T_6 = _GEN_197 & _warp_bar_exp_T_5; // @[warp_schedule.scala 98:54]
  wire [3:0] _warp_bar_belong_T_3 = ~_warp_bar_belong_T; // @[warp_schedule.scala 99:63]
  wire [3:0] _GEN_65 = 2'h1 == end_wg_id ? warp_bar_belong_1 : warp_bar_belong_0; // @[warp_schedule.scala 99:{60,60}]
  wire [3:0] _GEN_66 = 2'h2 == end_wg_id ? warp_bar_belong_2 : _GEN_65; // @[warp_schedule.scala 99:{60,60}]
  wire [3:0] _GEN_67 = 2'h3 == end_wg_id ? warp_bar_belong_3 : _GEN_66; // @[warp_schedule.scala 99:{60,60}]
  wire [3:0] _warp_bar_belong_T_4 = _GEN_67 & _warp_bar_belong_T_3; // @[warp_schedule.scala 99:60]
  wire [3:0] _GEN_81 = 2'h1 == end_wg_id ? warp_bar_cur_1 : warp_bar_cur_0; // @[warp_schedule.scala 103:{54,54}]
  wire [3:0] _GEN_82 = 2'h2 == end_wg_id ? warp_bar_cur_2 : _GEN_81; // @[warp_schedule.scala 103:{54,54}]
  wire [3:0] _GEN_83 = 2'h3 == end_wg_id ? warp_bar_cur_3 : _GEN_82; // @[warp_schedule.scala 103:{54,54}]
  wire [7:0] _GEN_198 = {{4'd0}, _GEN_83}; // @[warp_schedule.scala 103:54]
  wire [7:0] _warp_bar_cur_T_1 = _GEN_198 | _warp_bar_exp_T_4; // @[warp_schedule.scala 103:54]
  wire [3:0] _GEN_84 = 2'h0 == end_wg_id ? _warp_bar_cur_T_1[3:0] : _GEN_52; // @[warp_schedule.scala 103:{28,28}]
  wire [3:0] _GEN_85 = 2'h1 == end_wg_id ? _warp_bar_cur_T_1[3:0] : _GEN_53; // @[warp_schedule.scala 103:{28,28}]
  wire [3:0] _GEN_86 = 2'h2 == end_wg_id ? _warp_bar_cur_T_1[3:0] : _GEN_54; // @[warp_schedule.scala 103:{28,28}]
  wire [3:0] _GEN_87 = 2'h3 == end_wg_id ? _warp_bar_cur_T_1[3:0] : _GEN_55; // @[warp_schedule.scala 103:{28,28}]
  wire [3:0] _warp_bar_data_T = 4'h1 << io_warp_control_bits_ctrl_wid; // @[warp_schedule.scala 104:40]
  wire [3:0] _warp_bar_data_T_1 = warp_bar_data | _warp_bar_data_T; // @[warp_schedule.scala 104:34]
  wire [3:0] _warp_bar_data_T_2 = ~_GEN_67; // @[warp_schedule.scala 107:39]
  wire [3:0] _warp_bar_data_T_3 = warp_bar_data & _warp_bar_data_T_2; // @[warp_schedule.scala 107:36]
  wire [3:0] _warp_active_T_3 = _T_4 ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _warp_active_T_4 = _warp_bar_belong_T & _warp_active_T_3; // @[warp_schedule.scala 118:67]
  wire [3:0] _warp_active_T_5 = warp_active | _warp_active_T_4; // @[warp_schedule.scala 118:29]
  wire [3:0] _warp_active_T_7 = warp_end ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _warp_active_T_9 = _warp_active_T_7 & _warp_bar_data_T; // @[warp_schedule.scala 118:132]
  wire [3:0] _warp_active_T_10 = ~_warp_active_T_9; // @[warp_schedule.scala 118:106]
  wire [3:0] _warp_active_T_11 = _warp_active_T_5 & _warp_active_T_10; // @[warp_schedule.scala 118:103]
  wire [3:0] _warp_ready_T = warp_bar_data | io_scoreboard_busy; // @[warp_schedule.scala 119:35]
  wire [3:0] _warp_ready_T_1 = _warp_ready_T | io_exe_busy; // @[warp_schedule.scala 119:56]
  wire [3:0] _warp_ready_T_2 = ~warp_active; // @[warp_schedule.scala 119:73]
  wire [3:0] _warp_ready_T_3 = _warp_ready_T_1 | _warp_ready_T_2; // @[warp_schedule.scala 119:70]
  wire  _GEN_110 = 2'h0 == io_pc_rsp_bits_warpid ? 1'h0 : _GEN_4; // @[warp_schedule.scala 138:{47,47}]
  wire  _GEN_111 = 2'h1 == io_pc_rsp_bits_warpid ? 1'h0 : _GEN_5; // @[warp_schedule.scala 138:{47,47}]
  wire  _GEN_112 = 2'h2 == io_pc_rsp_bits_warpid ? 1'h0 : _GEN_6; // @[warp_schedule.scala 138:{47,47}]
  wire  _GEN_113 = 2'h3 == io_pc_rsp_bits_warpid ? 1'h0 : _GEN_7; // @[warp_schedule.scala 138:{47,47}]
  wire [1:0] _GEN_114 = 2'h0 == io_pc_rsp_bits_warpid ? 2'h1 : _GEN_8; // @[warp_schedule.scala 139:{44,44}]
  wire [1:0] _GEN_115 = 2'h1 == io_pc_rsp_bits_warpid ? 2'h1 : _GEN_9; // @[warp_schedule.scala 139:{44,44}]
  wire [1:0] _GEN_116 = 2'h2 == io_pc_rsp_bits_warpid ? 2'h1 : _GEN_10; // @[warp_schedule.scala 139:{44,44}]
  wire [1:0] _GEN_117 = 2'h3 == io_pc_rsp_bits_warpid ? 2'h1 : _GEN_11; // @[warp_schedule.scala 139:{44,44}]
  wire [31:0] _GEN_118 = 2'h0 == io_pc_rsp_bits_warpid ? io_pc_rsp_bits_addr : io_branch_bits_new_pc; // @[warp_schedule.scala 140:{44,44} 58:15]
  wire [31:0] _GEN_119 = 2'h1 == io_pc_rsp_bits_warpid ? io_pc_rsp_bits_addr : io_branch_bits_new_pc; // @[warp_schedule.scala 140:{44,44} 58:15]
  wire [31:0] _GEN_120 = 2'h2 == io_pc_rsp_bits_warpid ? io_pc_rsp_bits_addr : io_branch_bits_new_pc; // @[warp_schedule.scala 140:{44,44} 58:15]
  wire [31:0] _GEN_121 = 2'h3 == io_pc_rsp_bits_warpid ? io_pc_rsp_bits_addr : io_branch_bits_new_pc; // @[warp_schedule.scala 140:{44,44} 58:15]
  wire  _GEN_122 = _io_flushCache_valid_T_1 ? _GEN_110 : _GEN_4; // @[warp_schedule.scala 137:49]
  wire  _GEN_123 = _io_flushCache_valid_T_1 ? _GEN_111 : _GEN_5; // @[warp_schedule.scala 137:49]
  wire  _GEN_124 = _io_flushCache_valid_T_1 ? _GEN_112 : _GEN_6; // @[warp_schedule.scala 137:49]
  wire  _GEN_125 = _io_flushCache_valid_T_1 ? _GEN_113 : _GEN_7; // @[warp_schedule.scala 137:49]
  wire [1:0] _GEN_126 = _io_flushCache_valid_T_1 ? _GEN_114 : _GEN_8; // @[warp_schedule.scala 137:49]
  wire [1:0] _GEN_127 = _io_flushCache_valid_T_1 ? _GEN_115 : _GEN_9; // @[warp_schedule.scala 137:49]
  wire [1:0] _GEN_128 = _io_flushCache_valid_T_1 ? _GEN_116 : _GEN_10; // @[warp_schedule.scala 137:49]
  wire [1:0] _GEN_129 = _io_flushCache_valid_T_1 ? _GEN_117 : _GEN_11; // @[warp_schedule.scala 137:49]
  wire [31:0] _GEN_130 = _io_flushCache_valid_T_1 ? _GEN_118 : io_branch_bits_new_pc; // @[warp_schedule.scala 137:49 58:15]
  wire [31:0] _GEN_131 = _io_flushCache_valid_T_1 ? _GEN_119 : io_branch_bits_new_pc; // @[warp_schedule.scala 137:49 58:15]
  wire [31:0] _GEN_132 = _io_flushCache_valid_T_1 ? _GEN_120 : io_branch_bits_new_pc; // @[warp_schedule.scala 137:49 58:15]
  wire [31:0] _GEN_133 = _io_flushCache_valid_T_1 ? _GEN_121 : io_branch_bits_new_pc; // @[warp_schedule.scala 137:49 58:15]
  wire  _GEN_134 = 2'h0 == io_branch_bits_wid ? 1'h0 : _GEN_122; // @[warp_schedule.scala 144:{44,44}]
  wire  _GEN_135 = 2'h1 == io_branch_bits_wid ? 1'h0 : _GEN_123; // @[warp_schedule.scala 144:{44,44}]
  wire  _GEN_136 = 2'h2 == io_branch_bits_wid ? 1'h0 : _GEN_124; // @[warp_schedule.scala 144:{44,44}]
  wire  _GEN_137 = 2'h3 == io_branch_bits_wid ? 1'h0 : _GEN_125; // @[warp_schedule.scala 144:{44,44}]
  wire [1:0] _GEN_138 = 2'h0 == io_branch_bits_wid ? 2'h1 : _GEN_126; // @[warp_schedule.scala 145:{41,41}]
  wire [1:0] _GEN_139 = 2'h1 == io_branch_bits_wid ? 2'h1 : _GEN_127; // @[warp_schedule.scala 145:{41,41}]
  wire [1:0] _GEN_140 = 2'h2 == io_branch_bits_wid ? 2'h1 : _GEN_128; // @[warp_schedule.scala 145:{41,41}]
  wire [1:0] _GEN_141 = 2'h3 == io_branch_bits_wid ? 2'h1 : _GEN_129; // @[warp_schedule.scala 145:{41,41}]
  wire [31:0] _GEN_142 = 2'h0 == io_branch_bits_wid ? io_branch_bits_new_pc : _GEN_130; // @[warp_schedule.scala 146:{41,41}]
  wire [31:0] _GEN_143 = 2'h1 == io_branch_bits_wid ? io_branch_bits_new_pc : _GEN_131; // @[warp_schedule.scala 146:{41,41}]
  wire [31:0] _GEN_144 = 2'h2 == io_branch_bits_wid ? io_branch_bits_new_pc : _GEN_132; // @[warp_schedule.scala 146:{41,41}]
  wire [31:0] _GEN_145 = 2'h3 == io_branch_bits_wid ? io_branch_bits_new_pc : _GEN_133; // @[warp_schedule.scala 146:{41,41}]
  wire  _GEN_146 = io_branch_bits_wid == next_warp ? 1'h0 : _GEN_3; // @[warp_schedule.scala 126:18 148:41 149:20]
  wire  _GEN_147 = _io_flush_valid_T_1 ? _GEN_134 : _GEN_122; // @[warp_schedule.scala 143:45]
  wire  _GEN_148 = _io_flush_valid_T_1 ? _GEN_135 : _GEN_123; // @[warp_schedule.scala 143:45]
  wire  _GEN_149 = _io_flush_valid_T_1 ? _GEN_136 : _GEN_124; // @[warp_schedule.scala 143:45]
  wire  _GEN_150 = _io_flush_valid_T_1 ? _GEN_137 : _GEN_125; // @[warp_schedule.scala 143:45]
  wire [1:0] _GEN_151 = _io_flush_valid_T_1 ? _GEN_138 : _GEN_126; // @[warp_schedule.scala 143:45]
  wire [1:0] _GEN_152 = _io_flush_valid_T_1 ? _GEN_139 : _GEN_127; // @[warp_schedule.scala 143:45]
  wire [1:0] _GEN_153 = _io_flush_valid_T_1 ? _GEN_140 : _GEN_128; // @[warp_schedule.scala 143:45]
  wire [1:0] _GEN_154 = _io_flush_valid_T_1 ? _GEN_141 : _GEN_129; // @[warp_schedule.scala 143:45]
  wire [31:0] _GEN_155 = _io_flush_valid_T_1 ? _GEN_142 : _GEN_130; // @[warp_schedule.scala 143:45]
  wire [31:0] _GEN_156 = _io_flush_valid_T_1 ? _GEN_143 : _GEN_131; // @[warp_schedule.scala 143:45]
  wire [31:0] _GEN_157 = _io_flush_valid_T_1 ? _GEN_144 : _GEN_132; // @[warp_schedule.scala 143:45]
  wire [31:0] _GEN_158 = _io_flush_valid_T_1 ? _GEN_145 : _GEN_133; // @[warp_schedule.scala 143:45]
  wire  _GEN_159 = _io_flush_valid_T_1 ? _GEN_146 : _GEN_3; // @[warp_schedule.scala 126:18 143:45]
  wire  _GEN_160 = 2'h0 == io_warpReq_bits_wid ? 1'h0 : _GEN_147; // @[warp_schedule.scala 154:{45,45}]
  wire  _GEN_161 = 2'h1 == io_warpReq_bits_wid ? 1'h0 : _GEN_148; // @[warp_schedule.scala 154:{45,45}]
  wire  _GEN_162 = 2'h2 == io_warpReq_bits_wid ? 1'h0 : _GEN_149; // @[warp_schedule.scala 154:{45,45}]
  wire  _GEN_163 = 2'h3 == io_warpReq_bits_wid ? 1'h0 : _GEN_150; // @[warp_schedule.scala 154:{45,45}]
  wire [1:0] _GEN_164 = 2'h0 == io_warpReq_bits_wid ? 2'h1 : _GEN_151; // @[warp_schedule.scala 155:{42,42}]
  wire [1:0] _GEN_165 = 2'h1 == io_warpReq_bits_wid ? 2'h1 : _GEN_152; // @[warp_schedule.scala 155:{42,42}]
  wire [1:0] _GEN_166 = 2'h2 == io_warpReq_bits_wid ? 2'h1 : _GEN_153; // @[warp_schedule.scala 155:{42,42}]
  wire [1:0] _GEN_167 = 2'h3 == io_warpReq_bits_wid ? 2'h1 : _GEN_154; // @[warp_schedule.scala 155:{42,42}]
  wire [31:0] _GEN_168 = 2'h0 == io_warpReq_bits_wid ? io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch : _GEN_155; // @[warp_schedule.scala 156:{42,42}]
  wire [31:0] _GEN_169 = 2'h1 == io_warpReq_bits_wid ? io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch : _GEN_156; // @[warp_schedule.scala 156:{42,42}]
  wire [31:0] _GEN_170 = 2'h2 == io_warpReq_bits_wid ? io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch : _GEN_157; // @[warp_schedule.scala 156:{42,42}]
  wire [31:0] _GEN_171 = 2'h3 == io_warpReq_bits_wid ? io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch : _GEN_158; // @[warp_schedule.scala 156:{42,42}]
  wire  _GEN_172 = _T_4 ? _GEN_160 : _GEN_147; // @[warp_schedule.scala 153:26]
  wire  _GEN_173 = _T_4 ? _GEN_161 : _GEN_148; // @[warp_schedule.scala 153:26]
  wire  _GEN_174 = _T_4 ? _GEN_162 : _GEN_149; // @[warp_schedule.scala 153:26]
  wire  _GEN_175 = _T_4 ? _GEN_163 : _GEN_150; // @[warp_schedule.scala 153:26]
  wire [1:0] _GEN_176 = _T_4 ? _GEN_164 : _GEN_151; // @[warp_schedule.scala 153:26]
  wire [1:0] _GEN_177 = _T_4 ? _GEN_165 : _GEN_152; // @[warp_schedule.scala 153:26]
  wire [1:0] _GEN_178 = _T_4 ? _GEN_166 : _GEN_153; // @[warp_schedule.scala 153:26]
  wire [1:0] _GEN_179 = _T_4 ? _GEN_167 : _GEN_154; // @[warp_schedule.scala 153:26]
  wire [31:0] _GEN_180 = _T_4 ? _GEN_168 : _GEN_155; // @[warp_schedule.scala 153:26]
  wire [31:0] _GEN_181 = _T_4 ? _GEN_169 : _GEN_156; // @[warp_schedule.scala 153:26]
  wire [31:0] _GEN_182 = _T_4 ? _GEN_170 : _GEN_157; // @[warp_schedule.scala 153:26]
  wire [31:0] _GEN_183 = _T_4 ? _GEN_171 : _GEN_158; // @[warp_schedule.scala 153:26]
  PCcontrol PCcontrol ( // @[warp_schedule.scala 50:50]
    .clock(PCcontrol_clock),
    .reset(PCcontrol_reset),
    .io_New_PC(PCcontrol_io_New_PC),
    .io_PC_replay(PCcontrol_io_PC_replay),
    .io_PC_src(PCcontrol_io_PC_src),
    .io_PC_next(PCcontrol_io_PC_next)
  );
  PCcontrol PCcontrol_1 ( // @[warp_schedule.scala 50:50]
    .clock(PCcontrol_1_clock),
    .reset(PCcontrol_1_reset),
    .io_New_PC(PCcontrol_1_io_New_PC),
    .io_PC_replay(PCcontrol_1_io_PC_replay),
    .io_PC_src(PCcontrol_1_io_PC_src),
    .io_PC_next(PCcontrol_1_io_PC_next)
  );
  PCcontrol PCcontrol_2 ( // @[warp_schedule.scala 50:50]
    .clock(PCcontrol_2_clock),
    .reset(PCcontrol_2_reset),
    .io_New_PC(PCcontrol_2_io_New_PC),
    .io_PC_replay(PCcontrol_2_io_PC_replay),
    .io_PC_src(PCcontrol_2_io_PC_src),
    .io_PC_next(PCcontrol_2_io_PC_next)
  );
  PCcontrol PCcontrol_3 ( // @[warp_schedule.scala 50:50]
    .clock(PCcontrol_3_clock),
    .reset(PCcontrol_3_reset),
    .io_New_PC(PCcontrol_3_io_New_PC),
    .io_PC_replay(PCcontrol_3_io_PC_replay),
    .io_PC_src(PCcontrol_3_io_PC_src),
    .io_PC_next(PCcontrol_3_io_PC_next)
  );
  assign io_warpReq_ready = 1'h1; // @[warp_schedule.scala 37:19]
  assign io_warpRsp_valid = _warp_end_T & io_warp_control_bits_ctrl_simt_stack_op; // @[warp_schedule.scala 31:38]
  assign io_warpRsp_bits_wid = io_warp_control_bits_ctrl_wid; // @[warp_schedule.scala 39:22]
  assign io_wg_id_lookup = io_warp_control_bits_ctrl_barrier ? io_warp_control_bits_ctrl_wid : 2'h0; // @[warp_schedule.scala 75:23]
  assign io_pc_req_valid = io_pc_reset ? 1'h0 : _GEN_159; // @[warp_schedule.scala 160:20 162:20]
  assign io_pc_req_bits_addr = 2'h3 == next_warp ? pcControl_3_PC_next : _GEN_14; // @[warp_schedule.scala 72:{22,22}]
  assign io_pc_req_bits_warpid = pc_ready_0 ? 2'h0 : _GEN_104; // @[warp_schedule.scala 124:{22,32}]
  assign io_branch_ready = ~io_flushCache_valid; // @[warp_schedule.scala 34:21]
  assign io_warp_control_ready = ~_io_warp_control_ready_T & _io_branch_ready_T; // @[warp_schedule.scala 35:45]
  assign io_warp_ready = ~_warp_ready_T_3; // @[warp_schedule.scala 119:19]
  assign io_flush_valid = _io_warp_control_ready_T & io_branch_bits_jump | warp_end; // @[warp_schedule.scala 45:58]
  assign io_flush_bits = _io_flush_valid_T_1 ? io_branch_bits_wid : io_warp_control_bits_ctrl_wid; // @[warp_schedule.scala 46:21]
  assign io_flushCache_valid = io_pc_rsp_valid & io_pc_rsp_bits_status[0]; // @[warp_schedule.scala 47:39]
  assign io_flushCache_bits = io_pc_rsp_bits_warpid; // @[warp_schedule.scala 48:21]
  assign io_CTA2csr_valid = io_warpReq_valid; // @[warp_schedule.scala 42:19]
  assign io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count = io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count; // @[warp_schedule.scala 41:18]
  assign io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch = io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[warp_schedule.scala 41:18]
  assign io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch = io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch
    ; // @[warp_schedule.scala 41:18]
  assign io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch = io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch
    ; // @[warp_schedule.scala 41:18]
  assign io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch = io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[warp_schedule.scala 41:18]
  assign io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch = io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[warp_schedule.scala 41:18]
  assign io_CTA2csr_bits_wid = io_warpReq_bits_wid; // @[warp_schedule.scala 41:18]
  assign PCcontrol_clock = clock;
  assign PCcontrol_reset = reset;
  assign PCcontrol_io_New_PC = io_pc_reset ? 32'h0 : _GEN_180; // @[warp_schedule.scala 160:20 161:70]
  assign PCcontrol_io_PC_replay = io_pc_reset ? 1'h0 : _GEN_172; // @[warp_schedule.scala 160:20 161:101]
  assign PCcontrol_io_PC_src = io_pc_reset ? 2'h1 : _GEN_176; // @[warp_schedule.scala 160:20 161:56]
  assign PCcontrol_1_clock = clock;
  assign PCcontrol_1_reset = reset;
  assign PCcontrol_1_io_New_PC = io_pc_reset ? 32'h0 : _GEN_181; // @[warp_schedule.scala 160:20 161:70]
  assign PCcontrol_1_io_PC_replay = io_pc_reset ? 1'h0 : _GEN_173; // @[warp_schedule.scala 160:20 161:101]
  assign PCcontrol_1_io_PC_src = io_pc_reset ? 2'h1 : _GEN_177; // @[warp_schedule.scala 160:20 161:56]
  assign PCcontrol_2_clock = clock;
  assign PCcontrol_2_reset = reset;
  assign PCcontrol_2_io_New_PC = io_pc_reset ? 32'h0 : _GEN_182; // @[warp_schedule.scala 160:20 161:70]
  assign PCcontrol_2_io_PC_replay = io_pc_reset ? 1'h0 : _GEN_174; // @[warp_schedule.scala 160:20 161:101]
  assign PCcontrol_2_io_PC_src = io_pc_reset ? 2'h1 : _GEN_178; // @[warp_schedule.scala 160:20 161:56]
  assign PCcontrol_3_clock = clock;
  assign PCcontrol_3_reset = reset;
  assign PCcontrol_3_io_New_PC = io_pc_reset ? 32'h0 : _GEN_183; // @[warp_schedule.scala 160:20 161:70]
  assign PCcontrol_3_io_PC_replay = io_pc_reset ? 1'h0 : _GEN_175; // @[warp_schedule.scala 160:20 161:101]
  assign PCcontrol_3_io_PC_src = io_pc_reset ? 2'h1 : _GEN_179; // @[warp_schedule.scala 160:20 161:56]
  always @(posedge clock) begin
    if (reset) begin // @[warp_schedule.scala 65:27]
      current_warp <= 2'h0; // @[warp_schedule.scala 65:27]
    end else if (pc_ready_0) begin // @[warp_schedule.scala 124:22]
      current_warp <= 2'h0; // @[warp_schedule.scala 124:32]
    end else if (pc_ready_1) begin // @[warp_schedule.scala 124:22]
      current_warp <= 2'h1; // @[warp_schedule.scala 124:32]
    end else if (pc_ready_2) begin // @[warp_schedule.scala 124:22]
      current_warp <= 2'h2; // @[warp_schedule.scala 124:32]
    end else begin
      current_warp <= _GEN_102;
    end
    if (reset) begin // @[warp_schedule.scala 113:26]
      warp_active <= 4'h0; // @[warp_schedule.scala 113:26]
    end else begin
      warp_active <= _warp_active_T_11; // @[warp_schedule.scala 118:14]
    end
    if (reset) begin // @[warp_schedule.scala 77:27]
      warp_bar_cur_0 <= 4'h0; // @[warp_schedule.scala 77:27]
    end else if (_warp_end_T & ~io_warp_control_bits_ctrl_simt_stack_op) begin // @[warp_schedule.scala 102:72]
      if (_warp_bar_cur_T_1 == _GEN_197) begin // @[warp_schedule.scala 105:90]
        if (2'h0 == end_wg_id) begin // @[warp_schedule.scala 106:30]
          warp_bar_cur_0 <= 4'h0; // @[warp_schedule.scala 106:30]
        end else begin
          warp_bar_cur_0 <= _GEN_84;
        end
      end else begin
        warp_bar_cur_0 <= _GEN_84;
      end
    end else begin
      warp_bar_cur_0 <= _GEN_52;
    end
    if (reset) begin // @[warp_schedule.scala 77:27]
      warp_bar_cur_1 <= 4'h0; // @[warp_schedule.scala 77:27]
    end else if (_warp_end_T & ~io_warp_control_bits_ctrl_simt_stack_op) begin // @[warp_schedule.scala 102:72]
      if (_warp_bar_cur_T_1 == _GEN_197) begin // @[warp_schedule.scala 105:90]
        if (2'h1 == end_wg_id) begin // @[warp_schedule.scala 106:30]
          warp_bar_cur_1 <= 4'h0; // @[warp_schedule.scala 106:30]
        end else begin
          warp_bar_cur_1 <= _GEN_85;
        end
      end else begin
        warp_bar_cur_1 <= _GEN_85;
      end
    end else begin
      warp_bar_cur_1 <= _GEN_53;
    end
    if (reset) begin // @[warp_schedule.scala 77:27]
      warp_bar_cur_2 <= 4'h0; // @[warp_schedule.scala 77:27]
    end else if (_warp_end_T & ~io_warp_control_bits_ctrl_simt_stack_op) begin // @[warp_schedule.scala 102:72]
      if (_warp_bar_cur_T_1 == _GEN_197) begin // @[warp_schedule.scala 105:90]
        if (2'h2 == end_wg_id) begin // @[warp_schedule.scala 106:30]
          warp_bar_cur_2 <= 4'h0; // @[warp_schedule.scala 106:30]
        end else begin
          warp_bar_cur_2 <= _GEN_86;
        end
      end else begin
        warp_bar_cur_2 <= _GEN_86;
      end
    end else begin
      warp_bar_cur_2 <= _GEN_54;
    end
    if (reset) begin // @[warp_schedule.scala 77:27]
      warp_bar_cur_3 <= 4'h0; // @[warp_schedule.scala 77:27]
    end else if (_warp_end_T & ~io_warp_control_bits_ctrl_simt_stack_op) begin // @[warp_schedule.scala 102:72]
      if (_warp_bar_cur_T_1 == _GEN_197) begin // @[warp_schedule.scala 105:90]
        if (2'h3 == end_wg_id) begin // @[warp_schedule.scala 106:30]
          warp_bar_cur_3 <= 4'h0; // @[warp_schedule.scala 106:30]
        end else begin
          warp_bar_cur_3 <= _GEN_87;
        end
      end else begin
        warp_bar_cur_3 <= _GEN_87;
      end
    end else begin
      warp_bar_cur_3 <= _GEN_55;
    end
    if (reset) begin // @[warp_schedule.scala 78:27]
      warp_bar_exp_0 <= 4'h0; // @[warp_schedule.scala 78:27]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h0 == end_wg_id) begin // @[warp_schedule.scala 98:28]
        warp_bar_exp_0 <= _warp_bar_exp_T_6[3:0]; // @[warp_schedule.scala 98:28]
      end else begin
        warp_bar_exp_0 <= _GEN_48;
      end
    end else begin
      warp_bar_exp_0 <= _GEN_48;
    end
    if (reset) begin // @[warp_schedule.scala 78:27]
      warp_bar_exp_1 <= 4'h0; // @[warp_schedule.scala 78:27]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h1 == end_wg_id) begin // @[warp_schedule.scala 98:28]
        warp_bar_exp_1 <= _warp_bar_exp_T_6[3:0]; // @[warp_schedule.scala 98:28]
      end else begin
        warp_bar_exp_1 <= _GEN_49;
      end
    end else begin
      warp_bar_exp_1 <= _GEN_49;
    end
    if (reset) begin // @[warp_schedule.scala 78:27]
      warp_bar_exp_2 <= 4'h0; // @[warp_schedule.scala 78:27]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h2 == end_wg_id) begin // @[warp_schedule.scala 98:28]
        warp_bar_exp_2 <= _warp_bar_exp_T_6[3:0]; // @[warp_schedule.scala 98:28]
      end else begin
        warp_bar_exp_2 <= _GEN_50;
      end
    end else begin
      warp_bar_exp_2 <= _GEN_50;
    end
    if (reset) begin // @[warp_schedule.scala 78:27]
      warp_bar_exp_3 <= 4'h0; // @[warp_schedule.scala 78:27]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h3 == end_wg_id) begin // @[warp_schedule.scala 98:28]
        warp_bar_exp_3 <= _warp_bar_exp_T_6[3:0]; // @[warp_schedule.scala 98:28]
      end else begin
        warp_bar_exp_3 <= _GEN_51;
      end
    end else begin
      warp_bar_exp_3 <= _GEN_51;
    end
    if (reset) begin // @[warp_schedule.scala 81:28]
      warp_bar_lock_0 <= 1'h0; // @[warp_schedule.scala 81:28]
    end else begin
      warp_bar_lock_0 <= |warp_bar_exp_0; // @[warp_schedule.scala 101:16]
    end
    if (reset) begin // @[warp_schedule.scala 81:28]
      warp_bar_lock_1 <= 1'h0; // @[warp_schedule.scala 81:28]
    end else begin
      warp_bar_lock_1 <= |warp_bar_exp_1; // @[warp_schedule.scala 101:16]
    end
    if (reset) begin // @[warp_schedule.scala 81:28]
      warp_bar_lock_2 <= 1'h0; // @[warp_schedule.scala 81:28]
    end else begin
      warp_bar_lock_2 <= |warp_bar_exp_2; // @[warp_schedule.scala 101:16]
    end
    if (reset) begin // @[warp_schedule.scala 81:28]
      warp_bar_lock_3 <= 1'h0; // @[warp_schedule.scala 81:28]
    end else begin
      warp_bar_lock_3 <= |warp_bar_exp_3; // @[warp_schedule.scala 101:16]
    end
    if (reset) begin // @[warp_schedule.scala 87:28]
      warp_bar_data <= 4'h0; // @[warp_schedule.scala 87:28]
    end else if (_warp_end_T & ~io_warp_control_bits_ctrl_simt_stack_op) begin // @[warp_schedule.scala 102:72]
      if (_warp_bar_cur_T_1 == _GEN_197) begin // @[warp_schedule.scala 105:90]
        warp_bar_data <= _warp_bar_data_T_3; // @[warp_schedule.scala 107:20]
      end else begin
        warp_bar_data <= _warp_bar_data_T_1; // @[warp_schedule.scala 104:18]
      end
    end
    if (reset) begin // @[warp_schedule.scala 88:30]
      warp_bar_belong_0 <= 4'h0; // @[warp_schedule.scala 88:30]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h0 == end_wg_id) begin // @[warp_schedule.scala 99:31]
        warp_bar_belong_0 <= _warp_bar_belong_T_4; // @[warp_schedule.scala 99:31]
      end else begin
        warp_bar_belong_0 <= _GEN_44;
      end
    end else begin
      warp_bar_belong_0 <= _GEN_44;
    end
    if (reset) begin // @[warp_schedule.scala 88:30]
      warp_bar_belong_1 <= 4'h0; // @[warp_schedule.scala 88:30]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h1 == end_wg_id) begin // @[warp_schedule.scala 99:31]
        warp_bar_belong_1 <= _warp_bar_belong_T_4; // @[warp_schedule.scala 99:31]
      end else begin
        warp_bar_belong_1 <= _GEN_45;
      end
    end else begin
      warp_bar_belong_1 <= _GEN_45;
    end
    if (reset) begin // @[warp_schedule.scala 88:30]
      warp_bar_belong_2 <= 4'h0; // @[warp_schedule.scala 88:30]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h2 == end_wg_id) begin // @[warp_schedule.scala 99:31]
        warp_bar_belong_2 <= _warp_bar_belong_T_4; // @[warp_schedule.scala 99:31]
      end else begin
        warp_bar_belong_2 <= _GEN_46;
      end
    end else begin
      warp_bar_belong_2 <= _GEN_46;
    end
    if (reset) begin // @[warp_schedule.scala 88:30]
      warp_bar_belong_3 <= 4'h0; // @[warp_schedule.scala 88:30]
    end else if (io_warpRsp_valid) begin // @[warp_schedule.scala 97:24]
      if (2'h3 == end_wg_id) begin // @[warp_schedule.scala 99:31]
        warp_bar_belong_3 <= _warp_bar_belong_T_4; // @[warp_schedule.scala 99:31]
      end else begin
        warp_bar_belong_3 <= _GEN_47;
      end
    end else begin
      warp_bar_belong_3 <= _GEN_47;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  current_warp = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  warp_active = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  warp_bar_cur_0 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  warp_bar_cur_1 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  warp_bar_cur_2 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  warp_bar_cur_3 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  warp_bar_exp_0 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  warp_bar_exp_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  warp_bar_exp_2 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  warp_bar_exp_3 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  warp_bar_lock_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  warp_bar_lock_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  warp_bar_lock_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  warp_bar_lock_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  warp_bar_data = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  warp_bar_belong_0 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  warp_bar_belong_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  warp_bar_belong_2 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  warp_bar_belong_3 = _RAND_18[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Control(
  input  [31:0] io_inst,
  input  [31:0] io_pc,
  input  [1:0]  io_wid,
  output [31:0] io_control_inst,
  output [1:0]  io_control_wid,
  output        io_control_fp,
  output [1:0]  io_control_branch,
  output        io_control_simt_stack,
  output        io_control_simt_stack_op,
  output        io_control_barrier,
  output [1:0]  io_control_csr,
  output        io_control_reverse,
  output [1:0]  io_control_sel_alu2,
  output [1:0]  io_control_sel_alu1,
  output        io_control_isvec,
  output [1:0]  io_control_sel_alu3,
  output        io_control_mask,
  output [2:0]  io_control_sel_imm,
  output        io_control_mem_unsigned,
  output [5:0]  io_control_alu_fn,
  output        io_control_mem,
  output [1:0]  io_control_mem_cmd,
  output [1:0]  io_control_mop,
  output [4:0]  io_control_reg_idx1,
  output [4:0]  io_control_reg_idx2,
  output [4:0]  io_control_reg_idx3,
  output [4:0]  io_control_reg_idxw,
  output        io_control_wfd,
  output        io_control_fence,
  output        io_control_sfu,
  output        io_control_readmask,
  output        io_control_writemask,
  output        io_control_wxd,
  output [31:0] io_control_pc
);
  wire [31:0] _ctrlsignals_T = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_1 = 32'h100b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_3 = 32'hb == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_5 = 32'h400b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_7 = 32'h600b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_9 = 32'h500b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_11 = 32'h700b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_13 = 32'h300b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_14 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_15 = 32'h200200b == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_17 = 32'h200b == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_19 = 32'h1063 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_21 = 32'h63 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_23 = 32'h4063 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_25 = 32'h6063 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_27 = 32'h5063 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_29 = 32'h7063 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_30 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_31 = 32'h6f == _ctrlsignals_T_30; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_33 = 32'h67 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_35 = 32'h17 == _ctrlsignals_T_30; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_37 = 32'h1073 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_39 = 32'h2073 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_41 = 32'h3073 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_43 = 32'h5073 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_45 = 32'h6073 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_47 = 32'h7073 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_49 = 32'hf == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_51 = 32'h2003 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_53 = 32'h1003 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_55 = 32'h3 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_57 = 32'h5003 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_59 = 32'h4003 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_61 = 32'h2023 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_63 = 32'h1023 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_65 = 32'h23 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_67 = 32'h37 == _ctrlsignals_T_30; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_69 = 32'h13 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_71 = 32'h2013 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_73 = 32'h3013 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_75 = 32'h7013 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_77 = 32'h6013 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_79 = 32'h4013 == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_81 = 32'h33 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_83 = 32'h40000033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_85 = 32'h2033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_87 = 32'h3033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_89 = 32'h7033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_91 = 32'h6033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_93 = 32'h4033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_95 = 32'h1033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_97 = 32'h5033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_99 = 32'h40005033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_100 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_101 = 32'h1013 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_103 = 32'h5013 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_105 = 32'h40005013 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_107 = 32'h1b == _ctrlsignals_T; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_109 = 32'h2000033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_111 = 32'h2001033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_113 = 32'h2002033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_115 = 32'h2003033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_117 = 32'h2004033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_119 = 32'h2005033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_121 = 32'h2006033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_123 = 32'h2007033 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_124 = io_inst & 32'h600007f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_125 = 32'h43 == _ctrlsignals_T_124; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_127 = 32'h47 == _ctrlsignals_T_124; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_129 = 32'h4b == _ctrlsignals_T_124; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_131 = 32'h4f == _ctrlsignals_T_124; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_132 = io_inst & 32'hfe00007f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_133 = 32'h53 == _ctrlsignals_T_132; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_135 = 32'h8000053 == _ctrlsignals_T_132; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_137 = 32'h10000053 == _ctrlsignals_T_132; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_139 = 32'h18000053 == _ctrlsignals_T_132; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_140 = io_inst & 32'hfff0007f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_141 = 32'h58000053 == _ctrlsignals_T_140; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_143 = 32'h20000053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_145 = 32'h20001053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_147 = 32'h20002053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_149 = 32'h28000053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_151 = 32'h28001053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_153 = 32'hc0000053 == _ctrlsignals_T_140; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_155 = 32'hc0100053 == _ctrlsignals_T_140; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_159 = 32'ha0002053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_161 = 32'ha0001053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_163 = 32'ha0000053 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_164 = io_inst & 32'hfff0707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_165 = 32'he0001053 == _ctrlsignals_T_164; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_167 = 32'hd0000053 == _ctrlsignals_T_140; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_169 = 32'hd0100053 == _ctrlsignals_T_140; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_170 = io_inst & 32'h1df0707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_171 = 32'h6007 == _ctrlsignals_T_170; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_172 = io_inst & 32'h1c00707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_173 = 32'h8006007 == _ctrlsignals_T_172; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_175 = 32'hc006007 == _ctrlsignals_T_172; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_177 = 32'h6027 == _ctrlsignals_T_170; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_179 = 32'h8006027 == _ctrlsignals_T_172; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_181 = 32'hc006027 == _ctrlsignals_T_172; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_183 = 32'h90001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_185 = 32'h90005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_187 = 32'ha0001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_189 = 32'ha0005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_191 = 32'ha4001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_193 = 32'ha4005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_195 = 32'ha8001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_197 = 32'ha8005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_199 = 32'hac001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_201 = 32'hac005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_203 = 32'hb0001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_205 = 32'hb0005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_207 = 32'hb4001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_209 = 32'hb4005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_211 = 32'hb8001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_213 = 32'hb8005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_215 = 32'hbc001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_217 = 32'hbc005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_219 = 32'h57 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_221 = 32'h4057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_223 = 32'h3057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_225 = 32'h1057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_227 = 32'h5057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_229 = 32'h8001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_231 = 32'h8005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_233 = 32'h9c005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_235 = 32'h8000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_237 = 32'h8004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_239 = 32'hc004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_241 = 32'hc003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_243 = 32'h10001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_245 = 32'h10005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_247 = 32'h18001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_249 = 32'h18005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_251 = 32'h24000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_253 = 32'h24004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_255 = 32'h24003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_257 = 32'h28000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_259 = 32'h28004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_261 = 32'h28003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_263 = 32'h2c000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_265 = 32'h2c004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_267 = 32'h2c003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_269 = 32'h60000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_271 = 32'h60004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_273 = 32'h60003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_275 = 32'h64000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_277 = 32'h64004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_279 = 32'h64003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_281 = 32'h60001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_283 = 32'h60005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_285 = 32'h70001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_287 = 32'h70005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_289 = 32'h64001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_291 = 32'h64005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_293 = 32'h68000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_295 = 32'h68004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_297 = 32'h6c000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_299 = 32'h6c004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_301 = 32'h6c001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_303 = 32'h6c005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_305 = 32'h74005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_307 = 32'h7c005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_309 = 32'h94000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_311 = 32'h94004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_313 = 32'h94003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_315 = 32'ha0000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_317 = 32'ha0004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_319 = 32'ha0003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_321 = 32'ha4000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_323 = 32'ha4004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_325 = 32'ha4003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_327 = 32'h70000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_329 = 32'h70003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_331 = 32'h70004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_333 = 32'h74000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_335 = 32'h74003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_337 = 32'h74004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_339 = 32'h78003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_341 = 32'h78004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_343 = 32'h7c003057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_345 = 32'h7c004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_347 = 32'h64002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_349 = 32'h68002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_351 = 32'h6c002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_353 = 32'h60002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_355 = 32'h70002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_357 = 32'h74002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_359 = 32'h78002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_361 = 32'h7c002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_362 = io_inst & 32'hfdfff07f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_363 = 32'h5008a057 == _ctrlsignals_T_362; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_365 = 32'h5c000057 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_367 = 32'h5c004057 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_369 = 32'h5c003057 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_371 = 32'h94002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_373 = 32'h94006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_375 = 32'h9c002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_377 = 32'h9c006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_379 = 32'h90002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_381 = 32'h90006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_383 = 32'h98002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_385 = 32'h98006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_387 = 32'hb4002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_389 = 32'hb4006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_391 = 32'hbc002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_393 = 32'hbc006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_395 = 32'ha4002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_397 = 32'ha4006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_399 = 32'hac002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_401 = 32'hac006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_403 = 32'h8c002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_405 = 32'h8c006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_407 = 32'h88002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_409 = 32'h88006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_411 = 32'h84002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_413 = 32'h84006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_415 = 32'h80002057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_417 = 32'h80006057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_419 = 32'h80001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_421 = 32'h80005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_423 = 32'h84005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_424 = io_inst & 32'hfc0ff07f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_425 = 32'h4c001057 == _ctrlsignals_T_424; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_427 = 32'h10000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_429 = 32'h18000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_431 = 32'h14000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_433 = 32'h1c000057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_435 = 32'h10004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_437 = 32'h18004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_439 = 32'h14004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_441 = 32'h1c004057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_443 = 32'h20001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_445 = 32'h20005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_447 = 32'h24001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_449 = 32'h24005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_451 = 32'h28001057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_453 = 32'h28005057 == _ctrlsignals_T_100; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_459 = 32'h48001057 == _ctrlsignals_T_424; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_461 = 32'h48009057 == _ctrlsignals_T_424; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_463 = 32'h48011057 == _ctrlsignals_T_424; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_465 = 32'h48019057 == _ctrlsignals_T_424; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_467 = 32'h4c081057 == _ctrlsignals_T_424; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_469 = 32'h5e000057 == _ctrlsignals_T_164; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_471 = 32'h5e005057 == _ctrlsignals_T_164; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_473 = 32'h5e003057 == _ctrlsignals_T_164; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_475 = 32'h5e004057 == _ctrlsignals_T_164; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_476 = io_inst & 32'hfe0ff07f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_477 = 32'h42002057 == _ctrlsignals_T_476; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_478 = io_inst & 32'h8000707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_479 = 32'h7057 == _ctrlsignals_T_478; // @[Lookup.scala 31:38]
  wire [31:0] _ctrlsignals_T_480 = io_inst & 32'hc000707f; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_481 = 32'hc0007057 == _ctrlsignals_T_480; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_483 = 32'h80007057 == _ctrlsignals_T_14; // @[Lookup.scala 31:38]
  wire  _ctrlsignals_T_487 = _ctrlsignals_T_477 ? 1'h0 : _ctrlsignals_T_479 | (_ctrlsignals_T_481 | _ctrlsignals_T_483); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_517 = _ctrlsignals_T_417 | (_ctrlsignals_T_419 | (_ctrlsignals_T_421 | (_ctrlsignals_T_423 | (
    _ctrlsignals_T_425 | (_ctrlsignals_T_427 | (_ctrlsignals_T_429 | (_ctrlsignals_T_431 | (_ctrlsignals_T_433 | (
    _ctrlsignals_T_435 | (_ctrlsignals_T_437 | (_ctrlsignals_T_439 | (_ctrlsignals_T_441 | (_ctrlsignals_T_443 | (
    _ctrlsignals_T_445 | (_ctrlsignals_T_447 | (_ctrlsignals_T_449 | (_ctrlsignals_T_451 | (_ctrlsignals_T_453 | (
    _ctrlsignals_T_443 | (_ctrlsignals_T_445 | (_ctrlsignals_T_459 | (_ctrlsignals_T_461 | (_ctrlsignals_T_463 | (
    _ctrlsignals_T_465 | (_ctrlsignals_T_467 | (_ctrlsignals_T_469 | (_ctrlsignals_T_471 | (_ctrlsignals_T_473 | (
    _ctrlsignals_T_475 | _ctrlsignals_T_487))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_547 = _ctrlsignals_T_357 | (_ctrlsignals_T_359 | (_ctrlsignals_T_361 | (_ctrlsignals_T_363 | (
    _ctrlsignals_T_365 | (_ctrlsignals_T_367 | (_ctrlsignals_T_369 | (_ctrlsignals_T_371 | (_ctrlsignals_T_373 | (
    _ctrlsignals_T_375 | (_ctrlsignals_T_377 | (_ctrlsignals_T_379 | (_ctrlsignals_T_381 | (_ctrlsignals_T_383 | (
    _ctrlsignals_T_385 | (_ctrlsignals_T_387 | (_ctrlsignals_T_389 | (_ctrlsignals_T_391 | (_ctrlsignals_T_393 | (
    _ctrlsignals_T_395 | (_ctrlsignals_T_397 | (_ctrlsignals_T_399 | (_ctrlsignals_T_401 | (_ctrlsignals_T_403 | (
    _ctrlsignals_T_405 | (_ctrlsignals_T_407 | (_ctrlsignals_T_409 | (_ctrlsignals_T_411 | (_ctrlsignals_T_413 | (
    _ctrlsignals_T_415 | _ctrlsignals_T_517))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_577 = _ctrlsignals_T_297 | (_ctrlsignals_T_299 | (_ctrlsignals_T_301 | (_ctrlsignals_T_303 | (
    _ctrlsignals_T_305 | (_ctrlsignals_T_307 | (_ctrlsignals_T_309 | (_ctrlsignals_T_311 | (_ctrlsignals_T_313 | (
    _ctrlsignals_T_315 | (_ctrlsignals_T_317 | (_ctrlsignals_T_319 | (_ctrlsignals_T_321 | (_ctrlsignals_T_323 | (
    _ctrlsignals_T_325 | (_ctrlsignals_T_327 | (_ctrlsignals_T_329 | (_ctrlsignals_T_331 | (_ctrlsignals_T_333 | (
    _ctrlsignals_T_335 | (_ctrlsignals_T_337 | (_ctrlsignals_T_339 | (_ctrlsignals_T_341 | (_ctrlsignals_T_343 | (
    _ctrlsignals_T_345 | (_ctrlsignals_T_347 | (_ctrlsignals_T_349 | (_ctrlsignals_T_351 | (_ctrlsignals_T_353 | (
    _ctrlsignals_T_355 | _ctrlsignals_T_547))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_607 = _ctrlsignals_T_237 | (_ctrlsignals_T_239 | (_ctrlsignals_T_241 | (_ctrlsignals_T_243 | (
    _ctrlsignals_T_245 | (_ctrlsignals_T_247 | (_ctrlsignals_T_249 | (_ctrlsignals_T_251 | (_ctrlsignals_T_253 | (
    _ctrlsignals_T_255 | (_ctrlsignals_T_257 | (_ctrlsignals_T_259 | (_ctrlsignals_T_261 | (_ctrlsignals_T_263 | (
    _ctrlsignals_T_265 | (_ctrlsignals_T_267 | (_ctrlsignals_T_269 | (_ctrlsignals_T_271 | (_ctrlsignals_T_273 | (
    _ctrlsignals_T_275 | (_ctrlsignals_T_277 | (_ctrlsignals_T_279 | (_ctrlsignals_T_281 | (_ctrlsignals_T_283 | (
    _ctrlsignals_T_285 | (_ctrlsignals_T_287 | (_ctrlsignals_T_289 | (_ctrlsignals_T_291 | (_ctrlsignals_T_293 | (
    _ctrlsignals_T_295 | _ctrlsignals_T_577))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_637 = _ctrlsignals_T_177 | (_ctrlsignals_T_179 | (_ctrlsignals_T_181 | (_ctrlsignals_T_183 | (
    _ctrlsignals_T_185 | (_ctrlsignals_T_187 | (_ctrlsignals_T_189 | (_ctrlsignals_T_191 | (_ctrlsignals_T_193 | (
    _ctrlsignals_T_195 | (_ctrlsignals_T_197 | (_ctrlsignals_T_199 | (_ctrlsignals_T_201 | (_ctrlsignals_T_203 | (
    _ctrlsignals_T_205 | (_ctrlsignals_T_207 | (_ctrlsignals_T_209 | (_ctrlsignals_T_211 | (_ctrlsignals_T_213 | (
    _ctrlsignals_T_215 | (_ctrlsignals_T_217 | (_ctrlsignals_T_219 | (_ctrlsignals_T_221 | (_ctrlsignals_T_223 | (
    _ctrlsignals_T_225 | (_ctrlsignals_T_227 | (_ctrlsignals_T_229 | (_ctrlsignals_T_231 | (_ctrlsignals_T_233 | (
    _ctrlsignals_T_235 | _ctrlsignals_T_607))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_641 = _ctrlsignals_T_169 ? 1'h0 : _ctrlsignals_T_171 | (_ctrlsignals_T_173 | (_ctrlsignals_T_175
     | _ctrlsignals_T_637)); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_642 = _ctrlsignals_T_167 ? 1'h0 : _ctrlsignals_T_641; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_643 = _ctrlsignals_T_165 ? 1'h0 : _ctrlsignals_T_642; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_644 = _ctrlsignals_T_163 ? 1'h0 : _ctrlsignals_T_643; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_645 = _ctrlsignals_T_161 ? 1'h0 : _ctrlsignals_T_644; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_646 = _ctrlsignals_T_159 ? 1'h0 : _ctrlsignals_T_645; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_647 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_646; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_648 = _ctrlsignals_T_155 ? 1'h0 : _ctrlsignals_T_647; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_649 = _ctrlsignals_T_153 ? 1'h0 : _ctrlsignals_T_648; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_650 = _ctrlsignals_T_151 ? 1'h0 : _ctrlsignals_T_649; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_651 = _ctrlsignals_T_149 ? 1'h0 : _ctrlsignals_T_650; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_652 = _ctrlsignals_T_147 ? 1'h0 : _ctrlsignals_T_651; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_653 = _ctrlsignals_T_145 ? 1'h0 : _ctrlsignals_T_652; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_654 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_653; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_655 = _ctrlsignals_T_141 ? 1'h0 : _ctrlsignals_T_654; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_656 = _ctrlsignals_T_139 ? 1'h0 : _ctrlsignals_T_655; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_657 = _ctrlsignals_T_137 ? 1'h0 : _ctrlsignals_T_656; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_658 = _ctrlsignals_T_135 ? 1'h0 : _ctrlsignals_T_657; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_659 = _ctrlsignals_T_133 ? 1'h0 : _ctrlsignals_T_658; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_660 = _ctrlsignals_T_131 ? 1'h0 : _ctrlsignals_T_659; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_661 = _ctrlsignals_T_129 ? 1'h0 : _ctrlsignals_T_660; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_662 = _ctrlsignals_T_127 ? 1'h0 : _ctrlsignals_T_661; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_663 = _ctrlsignals_T_125 ? 1'h0 : _ctrlsignals_T_662; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_664 = _ctrlsignals_T_123 ? 1'h0 : _ctrlsignals_T_663; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_665 = _ctrlsignals_T_121 ? 1'h0 : _ctrlsignals_T_664; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_666 = _ctrlsignals_T_119 ? 1'h0 : _ctrlsignals_T_665; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_667 = _ctrlsignals_T_117 ? 1'h0 : _ctrlsignals_T_666; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_668 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_667; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_669 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_668; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_670 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_669; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_671 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_670; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_672 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_671; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_673 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_672; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_674 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_673; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_675 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_674; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_676 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_675; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_677 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_676; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_678 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_677; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_679 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_678; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_680 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_679; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_681 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_680; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_682 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_681; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_683 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_682; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_684 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_683; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_685 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_684; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_686 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_685; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_687 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_686; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_688 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_687; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_689 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_688; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_690 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_689; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_691 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_690; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_692 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_691; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_693 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_692; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_694 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_693; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_695 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_694; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_696 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_695; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_697 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_696; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_698 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_697; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_699 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_698; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_700 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_699; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_701 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_700; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_702 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_701; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_703 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_702; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_704 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_703; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_705 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_704; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_706 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_705; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_707 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_706; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_708 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_707; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_709 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_708; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_710 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_709; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_711 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_710; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_712 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_711; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_713 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_712; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_714 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_713; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_715 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_714; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_716 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_715; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_717 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_716; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_718 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_717; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_746 = _ctrlsignals_T_441 ? 1'h0 : _ctrlsignals_T_443 | (_ctrlsignals_T_445 | (_ctrlsignals_T_447
     | (_ctrlsignals_T_449 | (_ctrlsignals_T_451 | (_ctrlsignals_T_453 | (_ctrlsignals_T_443 | (_ctrlsignals_T_445 | (
    _ctrlsignals_T_459 | (_ctrlsignals_T_461 | (_ctrlsignals_T_463 | (_ctrlsignals_T_465 | _ctrlsignals_T_467)))))))))))
    ; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_747 = _ctrlsignals_T_439 ? 1'h0 : _ctrlsignals_T_746; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_748 = _ctrlsignals_T_437 ? 1'h0 : _ctrlsignals_T_747; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_749 = _ctrlsignals_T_435 ? 1'h0 : _ctrlsignals_T_748; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_750 = _ctrlsignals_T_433 ? 1'h0 : _ctrlsignals_T_749; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_751 = _ctrlsignals_T_431 ? 1'h0 : _ctrlsignals_T_750; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_752 = _ctrlsignals_T_429 ? 1'h0 : _ctrlsignals_T_751; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_753 = _ctrlsignals_T_427 ? 1'h0 : _ctrlsignals_T_752; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_758 = _ctrlsignals_T_417 ? 1'h0 : _ctrlsignals_T_419 | (_ctrlsignals_T_421 | (_ctrlsignals_T_423
     | (_ctrlsignals_T_425 | _ctrlsignals_T_753))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_759 = _ctrlsignals_T_415 ? 1'h0 : _ctrlsignals_T_758; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_760 = _ctrlsignals_T_413 ? 1'h0 : _ctrlsignals_T_759; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_761 = _ctrlsignals_T_411 ? 1'h0 : _ctrlsignals_T_760; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_762 = _ctrlsignals_T_409 ? 1'h0 : _ctrlsignals_T_761; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_763 = _ctrlsignals_T_407 ? 1'h0 : _ctrlsignals_T_762; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_764 = _ctrlsignals_T_405 ? 1'h0 : _ctrlsignals_T_763; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_765 = _ctrlsignals_T_403 ? 1'h0 : _ctrlsignals_T_764; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_766 = _ctrlsignals_T_401 ? 1'h0 : _ctrlsignals_T_765; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_767 = _ctrlsignals_T_399 ? 1'h0 : _ctrlsignals_T_766; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_768 = _ctrlsignals_T_397 ? 1'h0 : _ctrlsignals_T_767; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_769 = _ctrlsignals_T_395 ? 1'h0 : _ctrlsignals_T_768; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_770 = _ctrlsignals_T_393 ? 1'h0 : _ctrlsignals_T_769; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_771 = _ctrlsignals_T_391 ? 1'h0 : _ctrlsignals_T_770; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_772 = _ctrlsignals_T_389 ? 1'h0 : _ctrlsignals_T_771; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_773 = _ctrlsignals_T_387 ? 1'h0 : _ctrlsignals_T_772; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_774 = _ctrlsignals_T_385 ? 1'h0 : _ctrlsignals_T_773; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_775 = _ctrlsignals_T_383 ? 1'h0 : _ctrlsignals_T_774; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_776 = _ctrlsignals_T_381 ? 1'h0 : _ctrlsignals_T_775; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_777 = _ctrlsignals_T_379 ? 1'h0 : _ctrlsignals_T_776; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_778 = _ctrlsignals_T_377 ? 1'h0 : _ctrlsignals_T_777; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_779 = _ctrlsignals_T_375 ? 1'h0 : _ctrlsignals_T_778; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_780 = _ctrlsignals_T_373 ? 1'h0 : _ctrlsignals_T_779; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_781 = _ctrlsignals_T_371 ? 1'h0 : _ctrlsignals_T_780; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_782 = _ctrlsignals_T_369 ? 1'h0 : _ctrlsignals_T_781; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_783 = _ctrlsignals_T_367 ? 1'h0 : _ctrlsignals_T_782; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_784 = _ctrlsignals_T_365 ? 1'h0 : _ctrlsignals_T_783; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_785 = _ctrlsignals_T_363 ? 1'h0 : _ctrlsignals_T_784; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_786 = _ctrlsignals_T_361 ? 1'h0 : _ctrlsignals_T_785; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_787 = _ctrlsignals_T_359 ? 1'h0 : _ctrlsignals_T_786; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_788 = _ctrlsignals_T_357 ? 1'h0 : _ctrlsignals_T_787; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_789 = _ctrlsignals_T_355 ? 1'h0 : _ctrlsignals_T_788; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_790 = _ctrlsignals_T_353 ? 1'h0 : _ctrlsignals_T_789; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_791 = _ctrlsignals_T_351 ? 1'h0 : _ctrlsignals_T_790; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_792 = _ctrlsignals_T_349 ? 1'h0 : _ctrlsignals_T_791; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_793 = _ctrlsignals_T_347 ? 1'h0 : _ctrlsignals_T_792; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_794 = _ctrlsignals_T_345 ? 1'h0 : _ctrlsignals_T_793; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_795 = _ctrlsignals_T_343 ? 1'h0 : _ctrlsignals_T_794; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_796 = _ctrlsignals_T_341 ? 1'h0 : _ctrlsignals_T_795; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_797 = _ctrlsignals_T_339 ? 1'h0 : _ctrlsignals_T_796; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_798 = _ctrlsignals_T_337 ? 1'h0 : _ctrlsignals_T_797; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_799 = _ctrlsignals_T_335 ? 1'h0 : _ctrlsignals_T_798; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_800 = _ctrlsignals_T_333 ? 1'h0 : _ctrlsignals_T_799; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_801 = _ctrlsignals_T_331 ? 1'h0 : _ctrlsignals_T_800; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_802 = _ctrlsignals_T_329 ? 1'h0 : _ctrlsignals_T_801; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_803 = _ctrlsignals_T_327 ? 1'h0 : _ctrlsignals_T_802; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_804 = _ctrlsignals_T_325 ? 1'h0 : _ctrlsignals_T_803; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_805 = _ctrlsignals_T_323 ? 1'h0 : _ctrlsignals_T_804; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_806 = _ctrlsignals_T_321 ? 1'h0 : _ctrlsignals_T_805; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_807 = _ctrlsignals_T_319 ? 1'h0 : _ctrlsignals_T_806; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_808 = _ctrlsignals_T_317 ? 1'h0 : _ctrlsignals_T_807; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_809 = _ctrlsignals_T_315 ? 1'h0 : _ctrlsignals_T_808; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_810 = _ctrlsignals_T_313 ? 1'h0 : _ctrlsignals_T_809; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_811 = _ctrlsignals_T_311 ? 1'h0 : _ctrlsignals_T_810; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_812 = _ctrlsignals_T_309 ? 1'h0 : _ctrlsignals_T_811; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_817 = _ctrlsignals_T_299 ? 1'h0 : _ctrlsignals_T_301 | (_ctrlsignals_T_303 | (_ctrlsignals_T_305
     | (_ctrlsignals_T_307 | _ctrlsignals_T_812))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_818 = _ctrlsignals_T_297 ? 1'h0 : _ctrlsignals_T_817; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_819 = _ctrlsignals_T_295 ? 1'h0 : _ctrlsignals_T_818; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_820 = _ctrlsignals_T_293 ? 1'h0 : _ctrlsignals_T_819; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_827 = _ctrlsignals_T_279 ? 1'h0 : _ctrlsignals_T_281 | (_ctrlsignals_T_283 | (_ctrlsignals_T_285
     | (_ctrlsignals_T_287 | (_ctrlsignals_T_289 | (_ctrlsignals_T_291 | _ctrlsignals_T_820))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_828 = _ctrlsignals_T_277 ? 1'h0 : _ctrlsignals_T_827; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_829 = _ctrlsignals_T_275 ? 1'h0 : _ctrlsignals_T_828; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_830 = _ctrlsignals_T_273 ? 1'h0 : _ctrlsignals_T_829; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_831 = _ctrlsignals_T_271 ? 1'h0 : _ctrlsignals_T_830; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_832 = _ctrlsignals_T_269 ? 1'h0 : _ctrlsignals_T_831; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_833 = _ctrlsignals_T_267 ? 1'h0 : _ctrlsignals_T_832; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_834 = _ctrlsignals_T_265 ? 1'h0 : _ctrlsignals_T_833; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_835 = _ctrlsignals_T_263 ? 1'h0 : _ctrlsignals_T_834; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_836 = _ctrlsignals_T_261 ? 1'h0 : _ctrlsignals_T_835; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_837 = _ctrlsignals_T_259 ? 1'h0 : _ctrlsignals_T_836; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_838 = _ctrlsignals_T_257 ? 1'h0 : _ctrlsignals_T_837; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_839 = _ctrlsignals_T_255 ? 1'h0 : _ctrlsignals_T_838; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_840 = _ctrlsignals_T_253 ? 1'h0 : _ctrlsignals_T_839; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_841 = _ctrlsignals_T_251 ? 1'h0 : _ctrlsignals_T_840; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_846 = _ctrlsignals_T_241 ? 1'h0 : _ctrlsignals_T_243 | (_ctrlsignals_T_245 | (_ctrlsignals_T_247
     | (_ctrlsignals_T_249 | _ctrlsignals_T_841))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_847 = _ctrlsignals_T_239 ? 1'h0 : _ctrlsignals_T_846; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_848 = _ctrlsignals_T_237 ? 1'h0 : _ctrlsignals_T_847; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_849 = _ctrlsignals_T_235 ? 1'h0 : _ctrlsignals_T_848; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_855 = _ctrlsignals_T_223 ? 1'h0 : _ctrlsignals_T_225 | (_ctrlsignals_T_227 | (_ctrlsignals_T_229
     | (_ctrlsignals_T_231 | (_ctrlsignals_T_233 | _ctrlsignals_T_849)))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_856 = _ctrlsignals_T_221 ? 1'h0 : _ctrlsignals_T_855; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_857 = _ctrlsignals_T_219 ? 1'h0 : _ctrlsignals_T_856; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_876 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_183 | (_ctrlsignals_T_185 | (_ctrlsignals_T_187
     | (_ctrlsignals_T_189 | (_ctrlsignals_T_191 | (_ctrlsignals_T_193 | (_ctrlsignals_T_195 | (_ctrlsignals_T_197 | (
    _ctrlsignals_T_199 | (_ctrlsignals_T_201 | (_ctrlsignals_T_203 | (_ctrlsignals_T_205 | (_ctrlsignals_T_207 | (
    _ctrlsignals_T_209 | (_ctrlsignals_T_211 | (_ctrlsignals_T_213 | (_ctrlsignals_T_215 | (_ctrlsignals_T_217 |
    _ctrlsignals_T_857))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_877 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_876; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_878 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_877; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_879 = _ctrlsignals_T_175 ? 1'h0 : _ctrlsignals_T_878; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_880 = _ctrlsignals_T_173 ? 1'h0 : _ctrlsignals_T_879; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_881 = _ctrlsignals_T_171 ? 1'h0 : _ctrlsignals_T_880; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_905 = _ctrlsignals_T_123 ? 1'h0 : _ctrlsignals_T_125 | (_ctrlsignals_T_127 | (_ctrlsignals_T_129
     | (_ctrlsignals_T_131 | (_ctrlsignals_T_133 | (_ctrlsignals_T_135 | (_ctrlsignals_T_137 | (_ctrlsignals_T_139 | (
    _ctrlsignals_T_141 | (_ctrlsignals_T_143 | (_ctrlsignals_T_145 | (_ctrlsignals_T_147 | (_ctrlsignals_T_149 | (
    _ctrlsignals_T_151 | (_ctrlsignals_T_153 | (_ctrlsignals_T_155 | (_ctrlsignals_T_143 | (_ctrlsignals_T_159 | (
    _ctrlsignals_T_161 | (_ctrlsignals_T_163 | (_ctrlsignals_T_165 | (_ctrlsignals_T_167 | (_ctrlsignals_T_169 |
    _ctrlsignals_T_881)))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_906 = _ctrlsignals_T_121 ? 1'h0 : _ctrlsignals_T_905; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_907 = _ctrlsignals_T_119 ? 1'h0 : _ctrlsignals_T_906; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_908 = _ctrlsignals_T_117 ? 1'h0 : _ctrlsignals_T_907; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_909 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_908; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_910 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_909; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_911 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_910; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_912 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_911; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_913 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_912; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_914 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_913; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_915 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_914; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_916 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_915; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_917 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_916; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_918 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_917; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_919 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_918; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_920 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_919; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_921 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_920; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_922 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_921; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_923 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_922; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_924 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_923; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_925 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_924; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_926 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_925; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_927 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_926; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_928 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_927; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_929 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_928; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_930 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_929; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_931 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_930; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_932 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_931; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_933 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_932; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_934 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_933; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_935 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_934; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_936 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_935; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_937 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_936; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_938 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_937; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_939 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_938; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_940 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_939; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_941 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_940; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_942 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_941; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_943 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_942; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_944 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_943; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_945 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_944; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_946 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_945; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_947 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_946; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_948 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_947; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_949 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_948; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_950 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_949; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_951 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_950; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_952 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_951; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_953 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_952; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_954 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_953; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_955 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_954; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_956 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_955; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_957 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_956; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_958 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_957; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_959 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_958; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_960 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_959; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_961 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_960; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_962 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_961; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_963 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_962; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_964 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_963; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_965 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_964; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1201 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_15 | _ctrlsignals_T_17; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1202 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_1201; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1203 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_1202; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1204 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_1203; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1205 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_1204; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1206 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_1205; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1432 = _ctrlsignals_T_33 ? 2'h3 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1433 = _ctrlsignals_T_31 ? 2'h2 : _ctrlsignals_T_1432; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1434 = _ctrlsignals_T_29 ? 2'h1 : _ctrlsignals_T_1433; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1435 = _ctrlsignals_T_27 ? 2'h1 : _ctrlsignals_T_1434; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1436 = _ctrlsignals_T_25 ? 2'h1 : _ctrlsignals_T_1435; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1437 = _ctrlsignals_T_23 ? 2'h1 : _ctrlsignals_T_1436; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1438 = _ctrlsignals_T_21 ? 2'h1 : _ctrlsignals_T_1437; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1439 = _ctrlsignals_T_19 ? 2'h1 : _ctrlsignals_T_1438; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1440 = _ctrlsignals_T_17 ? 2'h0 : _ctrlsignals_T_1439; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1441 = _ctrlsignals_T_15 ? 2'h0 : _ctrlsignals_T_1440; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1442 = _ctrlsignals_T_13 ? 2'h1 : _ctrlsignals_T_1441; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1443 = _ctrlsignals_T_11 ? 2'h1 : _ctrlsignals_T_1442; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1444 = _ctrlsignals_T_9 ? 2'h1 : _ctrlsignals_T_1443; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1445 = _ctrlsignals_T_7 ? 2'h1 : _ctrlsignals_T_1444; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1446 = _ctrlsignals_T_5 ? 2'h1 : _ctrlsignals_T_1445; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1447 = _ctrlsignals_T_3 ? 2'h1 : _ctrlsignals_T_1446; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1923 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_17; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1925 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_13 | _ctrlsignals_T_1923; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1926 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_1925; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1927 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_1926; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1928 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_1927; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_1929 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_1928; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1930 = _ctrlsignals_T_483 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1931 = _ctrlsignals_T_481 ? 2'h2 : _ctrlsignals_T_1930; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1932 = _ctrlsignals_T_479 ? 2'h2 : _ctrlsignals_T_1931; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1933 = _ctrlsignals_T_477 ? 2'h0 : _ctrlsignals_T_1932; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1934 = _ctrlsignals_T_475 ? 2'h0 : _ctrlsignals_T_1933; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1935 = _ctrlsignals_T_473 ? 2'h0 : _ctrlsignals_T_1934; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1936 = _ctrlsignals_T_471 ? 2'h0 : _ctrlsignals_T_1935; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1937 = _ctrlsignals_T_469 ? 2'h0 : _ctrlsignals_T_1936; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1938 = _ctrlsignals_T_467 ? 2'h0 : _ctrlsignals_T_1937; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1939 = _ctrlsignals_T_465 ? 2'h0 : _ctrlsignals_T_1938; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1940 = _ctrlsignals_T_463 ? 2'h0 : _ctrlsignals_T_1939; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1941 = _ctrlsignals_T_461 ? 2'h0 : _ctrlsignals_T_1940; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1942 = _ctrlsignals_T_459 ? 2'h0 : _ctrlsignals_T_1941; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1943 = _ctrlsignals_T_445 ? 2'h0 : _ctrlsignals_T_1942; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1944 = _ctrlsignals_T_443 ? 2'h0 : _ctrlsignals_T_1943; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1945 = _ctrlsignals_T_453 ? 2'h0 : _ctrlsignals_T_1944; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1946 = _ctrlsignals_T_451 ? 2'h0 : _ctrlsignals_T_1945; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1947 = _ctrlsignals_T_449 ? 2'h0 : _ctrlsignals_T_1946; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1948 = _ctrlsignals_T_447 ? 2'h0 : _ctrlsignals_T_1947; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1949 = _ctrlsignals_T_445 ? 2'h0 : _ctrlsignals_T_1948; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1950 = _ctrlsignals_T_443 ? 2'h0 : _ctrlsignals_T_1949; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1951 = _ctrlsignals_T_441 ? 2'h0 : _ctrlsignals_T_1950; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1952 = _ctrlsignals_T_439 ? 2'h0 : _ctrlsignals_T_1951; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1953 = _ctrlsignals_T_437 ? 2'h0 : _ctrlsignals_T_1952; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1954 = _ctrlsignals_T_435 ? 2'h0 : _ctrlsignals_T_1953; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1955 = _ctrlsignals_T_433 ? 2'h0 : _ctrlsignals_T_1954; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1956 = _ctrlsignals_T_431 ? 2'h0 : _ctrlsignals_T_1955; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1957 = _ctrlsignals_T_429 ? 2'h0 : _ctrlsignals_T_1956; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1958 = _ctrlsignals_T_427 ? 2'h0 : _ctrlsignals_T_1957; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1959 = _ctrlsignals_T_425 ? 2'h0 : _ctrlsignals_T_1958; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1960 = _ctrlsignals_T_423 ? 2'h0 : _ctrlsignals_T_1959; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1961 = _ctrlsignals_T_421 ? 2'h0 : _ctrlsignals_T_1960; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1962 = _ctrlsignals_T_419 ? 2'h0 : _ctrlsignals_T_1961; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1963 = _ctrlsignals_T_417 ? 2'h0 : _ctrlsignals_T_1962; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1964 = _ctrlsignals_T_415 ? 2'h0 : _ctrlsignals_T_1963; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1965 = _ctrlsignals_T_413 ? 2'h0 : _ctrlsignals_T_1964; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1966 = _ctrlsignals_T_411 ? 2'h0 : _ctrlsignals_T_1965; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1967 = _ctrlsignals_T_409 ? 2'h0 : _ctrlsignals_T_1966; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1968 = _ctrlsignals_T_407 ? 2'h0 : _ctrlsignals_T_1967; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1969 = _ctrlsignals_T_405 ? 2'h0 : _ctrlsignals_T_1968; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1970 = _ctrlsignals_T_403 ? 2'h0 : _ctrlsignals_T_1969; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1971 = _ctrlsignals_T_401 ? 2'h0 : _ctrlsignals_T_1970; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1972 = _ctrlsignals_T_399 ? 2'h0 : _ctrlsignals_T_1971; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1973 = _ctrlsignals_T_397 ? 2'h0 : _ctrlsignals_T_1972; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1974 = _ctrlsignals_T_395 ? 2'h0 : _ctrlsignals_T_1973; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1975 = _ctrlsignals_T_393 ? 2'h0 : _ctrlsignals_T_1974; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1976 = _ctrlsignals_T_391 ? 2'h0 : _ctrlsignals_T_1975; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1977 = _ctrlsignals_T_389 ? 2'h0 : _ctrlsignals_T_1976; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1978 = _ctrlsignals_T_387 ? 2'h0 : _ctrlsignals_T_1977; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1979 = _ctrlsignals_T_385 ? 2'h0 : _ctrlsignals_T_1978; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1980 = _ctrlsignals_T_383 ? 2'h0 : _ctrlsignals_T_1979; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1981 = _ctrlsignals_T_381 ? 2'h0 : _ctrlsignals_T_1980; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1982 = _ctrlsignals_T_379 ? 2'h0 : _ctrlsignals_T_1981; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1983 = _ctrlsignals_T_377 ? 2'h0 : _ctrlsignals_T_1982; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1984 = _ctrlsignals_T_375 ? 2'h0 : _ctrlsignals_T_1983; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1985 = _ctrlsignals_T_373 ? 2'h0 : _ctrlsignals_T_1984; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1986 = _ctrlsignals_T_371 ? 2'h0 : _ctrlsignals_T_1985; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1987 = _ctrlsignals_T_369 ? 2'h0 : _ctrlsignals_T_1986; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1988 = _ctrlsignals_T_367 ? 2'h0 : _ctrlsignals_T_1987; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1989 = _ctrlsignals_T_365 ? 2'h0 : _ctrlsignals_T_1988; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1990 = _ctrlsignals_T_363 ? 2'h0 : _ctrlsignals_T_1989; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1991 = _ctrlsignals_T_361 ? 2'h0 : _ctrlsignals_T_1990; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1992 = _ctrlsignals_T_359 ? 2'h0 : _ctrlsignals_T_1991; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1993 = _ctrlsignals_T_357 ? 2'h0 : _ctrlsignals_T_1992; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1994 = _ctrlsignals_T_355 ? 2'h0 : _ctrlsignals_T_1993; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1995 = _ctrlsignals_T_353 ? 2'h0 : _ctrlsignals_T_1994; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1996 = _ctrlsignals_T_351 ? 2'h0 : _ctrlsignals_T_1995; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1997 = _ctrlsignals_T_349 ? 2'h0 : _ctrlsignals_T_1996; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1998 = _ctrlsignals_T_347 ? 2'h0 : _ctrlsignals_T_1997; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_1999 = _ctrlsignals_T_345 ? 2'h0 : _ctrlsignals_T_1998; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2000 = _ctrlsignals_T_343 ? 2'h0 : _ctrlsignals_T_1999; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2001 = _ctrlsignals_T_341 ? 2'h0 : _ctrlsignals_T_2000; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2002 = _ctrlsignals_T_339 ? 2'h0 : _ctrlsignals_T_2001; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2003 = _ctrlsignals_T_337 ? 2'h0 : _ctrlsignals_T_2002; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2004 = _ctrlsignals_T_335 ? 2'h0 : _ctrlsignals_T_2003; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2005 = _ctrlsignals_T_333 ? 2'h0 : _ctrlsignals_T_2004; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2006 = _ctrlsignals_T_331 ? 2'h0 : _ctrlsignals_T_2005; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2007 = _ctrlsignals_T_329 ? 2'h0 : _ctrlsignals_T_2006; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2008 = _ctrlsignals_T_327 ? 2'h0 : _ctrlsignals_T_2007; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2009 = _ctrlsignals_T_325 ? 2'h0 : _ctrlsignals_T_2008; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2010 = _ctrlsignals_T_323 ? 2'h0 : _ctrlsignals_T_2009; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2011 = _ctrlsignals_T_321 ? 2'h0 : _ctrlsignals_T_2010; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2012 = _ctrlsignals_T_319 ? 2'h0 : _ctrlsignals_T_2011; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2013 = _ctrlsignals_T_317 ? 2'h0 : _ctrlsignals_T_2012; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2014 = _ctrlsignals_T_315 ? 2'h0 : _ctrlsignals_T_2013; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2015 = _ctrlsignals_T_313 ? 2'h0 : _ctrlsignals_T_2014; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2016 = _ctrlsignals_T_311 ? 2'h0 : _ctrlsignals_T_2015; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2017 = _ctrlsignals_T_309 ? 2'h0 : _ctrlsignals_T_2016; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2018 = _ctrlsignals_T_307 ? 2'h0 : _ctrlsignals_T_2017; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2019 = _ctrlsignals_T_305 ? 2'h0 : _ctrlsignals_T_2018; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2020 = _ctrlsignals_T_303 ? 2'h0 : _ctrlsignals_T_2019; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2021 = _ctrlsignals_T_301 ? 2'h0 : _ctrlsignals_T_2020; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2022 = _ctrlsignals_T_299 ? 2'h0 : _ctrlsignals_T_2021; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2023 = _ctrlsignals_T_297 ? 2'h0 : _ctrlsignals_T_2022; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2024 = _ctrlsignals_T_295 ? 2'h0 : _ctrlsignals_T_2023; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2025 = _ctrlsignals_T_293 ? 2'h0 : _ctrlsignals_T_2024; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2026 = _ctrlsignals_T_291 ? 2'h0 : _ctrlsignals_T_2025; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2027 = _ctrlsignals_T_289 ? 2'h0 : _ctrlsignals_T_2026; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2028 = _ctrlsignals_T_287 ? 2'h0 : _ctrlsignals_T_2027; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2029 = _ctrlsignals_T_285 ? 2'h0 : _ctrlsignals_T_2028; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2030 = _ctrlsignals_T_283 ? 2'h0 : _ctrlsignals_T_2029; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2031 = _ctrlsignals_T_281 ? 2'h0 : _ctrlsignals_T_2030; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2032 = _ctrlsignals_T_279 ? 2'h0 : _ctrlsignals_T_2031; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2033 = _ctrlsignals_T_277 ? 2'h0 : _ctrlsignals_T_2032; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2034 = _ctrlsignals_T_275 ? 2'h0 : _ctrlsignals_T_2033; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2035 = _ctrlsignals_T_273 ? 2'h0 : _ctrlsignals_T_2034; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2036 = _ctrlsignals_T_271 ? 2'h0 : _ctrlsignals_T_2035; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2037 = _ctrlsignals_T_269 ? 2'h0 : _ctrlsignals_T_2036; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2038 = _ctrlsignals_T_267 ? 2'h0 : _ctrlsignals_T_2037; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2039 = _ctrlsignals_T_265 ? 2'h0 : _ctrlsignals_T_2038; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2040 = _ctrlsignals_T_263 ? 2'h0 : _ctrlsignals_T_2039; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2041 = _ctrlsignals_T_261 ? 2'h0 : _ctrlsignals_T_2040; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2042 = _ctrlsignals_T_259 ? 2'h0 : _ctrlsignals_T_2041; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2043 = _ctrlsignals_T_257 ? 2'h0 : _ctrlsignals_T_2042; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2044 = _ctrlsignals_T_255 ? 2'h0 : _ctrlsignals_T_2043; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2045 = _ctrlsignals_T_253 ? 2'h0 : _ctrlsignals_T_2044; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2046 = _ctrlsignals_T_251 ? 2'h0 : _ctrlsignals_T_2045; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2047 = _ctrlsignals_T_249 ? 2'h0 : _ctrlsignals_T_2046; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2048 = _ctrlsignals_T_247 ? 2'h0 : _ctrlsignals_T_2047; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2049 = _ctrlsignals_T_245 ? 2'h0 : _ctrlsignals_T_2048; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2050 = _ctrlsignals_T_243 ? 2'h0 : _ctrlsignals_T_2049; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2051 = _ctrlsignals_T_241 ? 2'h0 : _ctrlsignals_T_2050; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2052 = _ctrlsignals_T_239 ? 2'h0 : _ctrlsignals_T_2051; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2053 = _ctrlsignals_T_237 ? 2'h0 : _ctrlsignals_T_2052; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2054 = _ctrlsignals_T_235 ? 2'h0 : _ctrlsignals_T_2053; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2055 = _ctrlsignals_T_233 ? 2'h0 : _ctrlsignals_T_2054; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2056 = _ctrlsignals_T_231 ? 2'h0 : _ctrlsignals_T_2055; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2057 = _ctrlsignals_T_229 ? 2'h0 : _ctrlsignals_T_2056; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2058 = _ctrlsignals_T_227 ? 2'h0 : _ctrlsignals_T_2057; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2059 = _ctrlsignals_T_225 ? 2'h0 : _ctrlsignals_T_2058; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2060 = _ctrlsignals_T_223 ? 2'h0 : _ctrlsignals_T_2059; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2061 = _ctrlsignals_T_221 ? 2'h0 : _ctrlsignals_T_2060; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2062 = _ctrlsignals_T_219 ? 2'h0 : _ctrlsignals_T_2061; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2063 = _ctrlsignals_T_217 ? 2'h0 : _ctrlsignals_T_2062; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2064 = _ctrlsignals_T_215 ? 2'h0 : _ctrlsignals_T_2063; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2065 = _ctrlsignals_T_213 ? 2'h0 : _ctrlsignals_T_2064; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2066 = _ctrlsignals_T_211 ? 2'h0 : _ctrlsignals_T_2065; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2067 = _ctrlsignals_T_209 ? 2'h0 : _ctrlsignals_T_2066; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2068 = _ctrlsignals_T_207 ? 2'h0 : _ctrlsignals_T_2067; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2069 = _ctrlsignals_T_205 ? 2'h0 : _ctrlsignals_T_2068; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2070 = _ctrlsignals_T_203 ? 2'h0 : _ctrlsignals_T_2069; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2071 = _ctrlsignals_T_201 ? 2'h0 : _ctrlsignals_T_2070; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2072 = _ctrlsignals_T_199 ? 2'h0 : _ctrlsignals_T_2071; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2073 = _ctrlsignals_T_197 ? 2'h0 : _ctrlsignals_T_2072; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2074 = _ctrlsignals_T_195 ? 2'h0 : _ctrlsignals_T_2073; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2075 = _ctrlsignals_T_193 ? 2'h0 : _ctrlsignals_T_2074; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2076 = _ctrlsignals_T_191 ? 2'h0 : _ctrlsignals_T_2075; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2077 = _ctrlsignals_T_189 ? 2'h0 : _ctrlsignals_T_2076; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2078 = _ctrlsignals_T_187 ? 2'h0 : _ctrlsignals_T_2077; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2079 = _ctrlsignals_T_185 ? 2'h0 : _ctrlsignals_T_2078; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2080 = _ctrlsignals_T_183 ? 2'h0 : _ctrlsignals_T_2079; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2081 = _ctrlsignals_T_181 ? 2'h0 : _ctrlsignals_T_2080; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2082 = _ctrlsignals_T_179 ? 2'h0 : _ctrlsignals_T_2081; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2083 = _ctrlsignals_T_177 ? 2'h0 : _ctrlsignals_T_2082; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2084 = _ctrlsignals_T_175 ? 2'h0 : _ctrlsignals_T_2083; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2085 = _ctrlsignals_T_173 ? 2'h0 : _ctrlsignals_T_2084; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2086 = _ctrlsignals_T_171 ? 2'h0 : _ctrlsignals_T_2085; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2087 = _ctrlsignals_T_169 ? 2'h0 : _ctrlsignals_T_2086; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2088 = _ctrlsignals_T_167 ? 2'h0 : _ctrlsignals_T_2087; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2089 = _ctrlsignals_T_165 ? 2'h0 : _ctrlsignals_T_2088; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2090 = _ctrlsignals_T_163 ? 2'h0 : _ctrlsignals_T_2089; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2091 = _ctrlsignals_T_161 ? 2'h0 : _ctrlsignals_T_2090; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2092 = _ctrlsignals_T_159 ? 2'h0 : _ctrlsignals_T_2091; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2093 = _ctrlsignals_T_143 ? 2'h0 : _ctrlsignals_T_2092; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2094 = _ctrlsignals_T_155 ? 2'h0 : _ctrlsignals_T_2093; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2095 = _ctrlsignals_T_153 ? 2'h0 : _ctrlsignals_T_2094; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2096 = _ctrlsignals_T_151 ? 2'h0 : _ctrlsignals_T_2095; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2097 = _ctrlsignals_T_149 ? 2'h0 : _ctrlsignals_T_2096; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2098 = _ctrlsignals_T_147 ? 2'h0 : _ctrlsignals_T_2097; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2099 = _ctrlsignals_T_145 ? 2'h0 : _ctrlsignals_T_2098; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2100 = _ctrlsignals_T_143 ? 2'h0 : _ctrlsignals_T_2099; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2101 = _ctrlsignals_T_141 ? 2'h0 : _ctrlsignals_T_2100; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2102 = _ctrlsignals_T_139 ? 2'h0 : _ctrlsignals_T_2101; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2103 = _ctrlsignals_T_137 ? 2'h0 : _ctrlsignals_T_2102; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2104 = _ctrlsignals_T_135 ? 2'h0 : _ctrlsignals_T_2103; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2105 = _ctrlsignals_T_133 ? 2'h0 : _ctrlsignals_T_2104; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2106 = _ctrlsignals_T_131 ? 2'h0 : _ctrlsignals_T_2105; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2107 = _ctrlsignals_T_129 ? 2'h0 : _ctrlsignals_T_2106; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2108 = _ctrlsignals_T_127 ? 2'h0 : _ctrlsignals_T_2107; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2109 = _ctrlsignals_T_125 ? 2'h0 : _ctrlsignals_T_2108; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2110 = _ctrlsignals_T_123 ? 2'h0 : _ctrlsignals_T_2109; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2111 = _ctrlsignals_T_121 ? 2'h0 : _ctrlsignals_T_2110; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2112 = _ctrlsignals_T_119 ? 2'h0 : _ctrlsignals_T_2111; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2113 = _ctrlsignals_T_117 ? 2'h0 : _ctrlsignals_T_2112; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2114 = _ctrlsignals_T_115 ? 2'h0 : _ctrlsignals_T_2113; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2115 = _ctrlsignals_T_113 ? 2'h0 : _ctrlsignals_T_2114; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2116 = _ctrlsignals_T_111 ? 2'h0 : _ctrlsignals_T_2115; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2117 = _ctrlsignals_T_109 ? 2'h0 : _ctrlsignals_T_2116; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2118 = _ctrlsignals_T_107 ? 2'h0 : _ctrlsignals_T_2117; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2119 = _ctrlsignals_T_105 ? 2'h0 : _ctrlsignals_T_2118; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2120 = _ctrlsignals_T_103 ? 2'h0 : _ctrlsignals_T_2119; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2121 = _ctrlsignals_T_101 ? 2'h0 : _ctrlsignals_T_2120; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2122 = _ctrlsignals_T_99 ? 2'h0 : _ctrlsignals_T_2121; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2123 = _ctrlsignals_T_97 ? 2'h0 : _ctrlsignals_T_2122; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2124 = _ctrlsignals_T_95 ? 2'h0 : _ctrlsignals_T_2123; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2125 = _ctrlsignals_T_93 ? 2'h0 : _ctrlsignals_T_2124; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2126 = _ctrlsignals_T_91 ? 2'h0 : _ctrlsignals_T_2125; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2127 = _ctrlsignals_T_89 ? 2'h0 : _ctrlsignals_T_2126; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2128 = _ctrlsignals_T_87 ? 2'h0 : _ctrlsignals_T_2127; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2129 = _ctrlsignals_T_85 ? 2'h0 : _ctrlsignals_T_2128; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2130 = _ctrlsignals_T_83 ? 2'h0 : _ctrlsignals_T_2129; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2131 = _ctrlsignals_T_81 ? 2'h0 : _ctrlsignals_T_2130; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2132 = _ctrlsignals_T_79 ? 2'h0 : _ctrlsignals_T_2131; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2133 = _ctrlsignals_T_77 ? 2'h0 : _ctrlsignals_T_2132; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2134 = _ctrlsignals_T_75 ? 2'h0 : _ctrlsignals_T_2133; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2135 = _ctrlsignals_T_73 ? 2'h0 : _ctrlsignals_T_2134; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2136 = _ctrlsignals_T_71 ? 2'h0 : _ctrlsignals_T_2135; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2137 = _ctrlsignals_T_69 ? 2'h0 : _ctrlsignals_T_2136; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2138 = _ctrlsignals_T_67 ? 2'h0 : _ctrlsignals_T_2137; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2139 = _ctrlsignals_T_65 ? 2'h0 : _ctrlsignals_T_2138; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2140 = _ctrlsignals_T_63 ? 2'h0 : _ctrlsignals_T_2139; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2141 = _ctrlsignals_T_61 ? 2'h0 : _ctrlsignals_T_2140; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2142 = _ctrlsignals_T_59 ? 2'h0 : _ctrlsignals_T_2141; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2143 = _ctrlsignals_T_57 ? 2'h0 : _ctrlsignals_T_2142; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2144 = _ctrlsignals_T_55 ? 2'h0 : _ctrlsignals_T_2143; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2145 = _ctrlsignals_T_53 ? 2'h0 : _ctrlsignals_T_2144; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2146 = _ctrlsignals_T_51 ? 2'h0 : _ctrlsignals_T_2145; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2147 = _ctrlsignals_T_49 ? 2'h0 : _ctrlsignals_T_2146; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2148 = _ctrlsignals_T_47 ? 2'h3 : _ctrlsignals_T_2147; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2149 = _ctrlsignals_T_45 ? 2'h2 : _ctrlsignals_T_2148; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2150 = _ctrlsignals_T_43 ? 2'h1 : _ctrlsignals_T_2149; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2151 = _ctrlsignals_T_41 ? 2'h3 : _ctrlsignals_T_2150; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2152 = _ctrlsignals_T_39 ? 2'h2 : _ctrlsignals_T_2151; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2153 = _ctrlsignals_T_37 ? 2'h1 : _ctrlsignals_T_2152; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2154 = _ctrlsignals_T_35 ? 2'h0 : _ctrlsignals_T_2153; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2155 = _ctrlsignals_T_33 ? 2'h0 : _ctrlsignals_T_2154; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2156 = _ctrlsignals_T_31 ? 2'h0 : _ctrlsignals_T_2155; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2157 = _ctrlsignals_T_29 ? 2'h0 : _ctrlsignals_T_2156; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2158 = _ctrlsignals_T_27 ? 2'h0 : _ctrlsignals_T_2157; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2159 = _ctrlsignals_T_25 ? 2'h0 : _ctrlsignals_T_2158; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2160 = _ctrlsignals_T_23 ? 2'h0 : _ctrlsignals_T_2159; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2161 = _ctrlsignals_T_21 ? 2'h0 : _ctrlsignals_T_2160; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2162 = _ctrlsignals_T_19 ? 2'h0 : _ctrlsignals_T_2161; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2163 = _ctrlsignals_T_17 ? 2'h0 : _ctrlsignals_T_2162; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2164 = _ctrlsignals_T_15 ? 2'h0 : _ctrlsignals_T_2163; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2165 = _ctrlsignals_T_13 ? 2'h0 : _ctrlsignals_T_2164; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2166 = _ctrlsignals_T_11 ? 2'h0 : _ctrlsignals_T_2165; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2167 = _ctrlsignals_T_9 ? 2'h0 : _ctrlsignals_T_2166; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2168 = _ctrlsignals_T_7 ? 2'h0 : _ctrlsignals_T_2167; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2169 = _ctrlsignals_T_5 ? 2'h0 : _ctrlsignals_T_2168; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2170 = _ctrlsignals_T_3 ? 2'h0 : _ctrlsignals_T_2169; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2201 = _ctrlsignals_T_423 ? 1'h0 : _ctrlsignals_T_425 | _ctrlsignals_T_753; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2228 = _ctrlsignals_T_369 ? 1'h0 : _ctrlsignals_T_371 | (_ctrlsignals_T_373 | (_ctrlsignals_T_375
     | (_ctrlsignals_T_377 | (_ctrlsignals_T_379 | (_ctrlsignals_T_381 | (_ctrlsignals_T_383 | (_ctrlsignals_T_385 | (
    _ctrlsignals_T_387 | (_ctrlsignals_T_389 | (_ctrlsignals_T_391 | (_ctrlsignals_T_393 | (_ctrlsignals_T_395 | (
    _ctrlsignals_T_397 | (_ctrlsignals_T_399 | (_ctrlsignals_T_401 | (_ctrlsignals_T_403 | (_ctrlsignals_T_405 | (
    _ctrlsignals_T_407 | (_ctrlsignals_T_409 | (_ctrlsignals_T_411 | (_ctrlsignals_T_413 | (_ctrlsignals_T_415 | (
    _ctrlsignals_T_417 | (_ctrlsignals_T_419 | (_ctrlsignals_T_421 | _ctrlsignals_T_2201))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2229 = _ctrlsignals_T_367 ? 1'h0 : _ctrlsignals_T_2228; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2230 = _ctrlsignals_T_365 ? 1'h0 : _ctrlsignals_T_2229; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2231 = _ctrlsignals_T_363 ? 1'h0 : _ctrlsignals_T_2230; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2232 = _ctrlsignals_T_361 ? 1'h0 : _ctrlsignals_T_2231; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2233 = _ctrlsignals_T_359 ? 1'h0 : _ctrlsignals_T_2232; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2234 = _ctrlsignals_T_357 ? 1'h0 : _ctrlsignals_T_2233; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2235 = _ctrlsignals_T_355 ? 1'h0 : _ctrlsignals_T_2234; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2236 = _ctrlsignals_T_353 ? 1'h0 : _ctrlsignals_T_2235; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2237 = _ctrlsignals_T_351 ? 1'h0 : _ctrlsignals_T_2236; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2238 = _ctrlsignals_T_349 ? 1'h0 : _ctrlsignals_T_2237; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2239 = _ctrlsignals_T_347 ? 1'h0 : _ctrlsignals_T_2238; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2240 = _ctrlsignals_T_345 ? 1'h0 : _ctrlsignals_T_2239; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2241 = _ctrlsignals_T_343 ? 1'h0 : _ctrlsignals_T_2240; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2242 = _ctrlsignals_T_341 ? 1'h0 : _ctrlsignals_T_2241; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2243 = _ctrlsignals_T_339 ? 1'h0 : _ctrlsignals_T_2242; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2244 = _ctrlsignals_T_337 ? 1'h0 : _ctrlsignals_T_2243; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2245 = _ctrlsignals_T_335 ? 1'h0 : _ctrlsignals_T_2244; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2246 = _ctrlsignals_T_333 ? 1'h0 : _ctrlsignals_T_2245; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2247 = _ctrlsignals_T_331 ? 1'h0 : _ctrlsignals_T_2246; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2248 = _ctrlsignals_T_329 ? 1'h0 : _ctrlsignals_T_2247; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2249 = _ctrlsignals_T_327 ? 1'h0 : _ctrlsignals_T_2248; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2259 = _ctrlsignals_T_307 ? 1'h0 : _ctrlsignals_T_309 | (_ctrlsignals_T_311 | (_ctrlsignals_T_313
     | (_ctrlsignals_T_315 | (_ctrlsignals_T_317 | (_ctrlsignals_T_319 | (_ctrlsignals_T_321 | (_ctrlsignals_T_323 | (
    _ctrlsignals_T_325 | _ctrlsignals_T_2249)))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2260 = _ctrlsignals_T_305 ? 1'h0 : _ctrlsignals_T_2259; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2269 = _ctrlsignals_T_287 ? 1'h0 : _ctrlsignals_T_289 | (_ctrlsignals_T_291 | (_ctrlsignals_T_293
     | (_ctrlsignals_T_295 | (_ctrlsignals_T_297 | (_ctrlsignals_T_299 | (_ctrlsignals_T_301 | (_ctrlsignals_T_303 |
    _ctrlsignals_T_2260))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2270 = _ctrlsignals_T_285 ? 1'h0 : _ctrlsignals_T_2269; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2271 = _ctrlsignals_T_283 ? 1'h0 : _ctrlsignals_T_2270; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2272 = _ctrlsignals_T_281 ? 1'h0 : _ctrlsignals_T_2271; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2273 = _ctrlsignals_T_279 ? 1'h0 : _ctrlsignals_T_2272; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2274 = _ctrlsignals_T_277 ? 1'h0 : _ctrlsignals_T_2273; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2275 = _ctrlsignals_T_275 ? 1'h0 : _ctrlsignals_T_2274; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2276 = _ctrlsignals_T_273 ? 1'h0 : _ctrlsignals_T_2275; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2277 = _ctrlsignals_T_271 ? 1'h0 : _ctrlsignals_T_2276; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2278 = _ctrlsignals_T_269 ? 1'h0 : _ctrlsignals_T_2277; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2279 = _ctrlsignals_T_267 ? 1'h0 : _ctrlsignals_T_2278; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2280 = _ctrlsignals_T_265 ? 1'h0 : _ctrlsignals_T_2279; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2281 = _ctrlsignals_T_263 ? 1'h0 : _ctrlsignals_T_2280; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2282 = _ctrlsignals_T_261 ? 1'h0 : _ctrlsignals_T_2281; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2283 = _ctrlsignals_T_259 ? 1'h0 : _ctrlsignals_T_2282; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2284 = _ctrlsignals_T_257 ? 1'h0 : _ctrlsignals_T_2283; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2285 = _ctrlsignals_T_255 ? 1'h0 : _ctrlsignals_T_2284; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2286 = _ctrlsignals_T_253 ? 1'h0 : _ctrlsignals_T_2285; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2287 = _ctrlsignals_T_251 ? 1'h0 : _ctrlsignals_T_2286; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2288 = _ctrlsignals_T_249 ? 1'h0 : _ctrlsignals_T_2287; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2289 = _ctrlsignals_T_247 ? 1'h0 : _ctrlsignals_T_2288; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2290 = _ctrlsignals_T_245 ? 1'h0 : _ctrlsignals_T_2289; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2291 = _ctrlsignals_T_243 ? 1'h0 : _ctrlsignals_T_2290; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2292 = _ctrlsignals_T_241 ? 1'h0 : _ctrlsignals_T_2291; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2293 = _ctrlsignals_T_239 ? 1'h0 : _ctrlsignals_T_2292; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2296 = _ctrlsignals_T_233 ? 1'h0 : _ctrlsignals_T_235 | (_ctrlsignals_T_237 | _ctrlsignals_T_2293
    ); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2312 = _ctrlsignals_T_201 ? 1'h0 : _ctrlsignals_T_203 | (_ctrlsignals_T_205 | (_ctrlsignals_T_207
     | (_ctrlsignals_T_209 | (_ctrlsignals_T_211 | (_ctrlsignals_T_213 | (_ctrlsignals_T_215 | (_ctrlsignals_T_217 | (
    _ctrlsignals_T_219 | (_ctrlsignals_T_221 | (_ctrlsignals_T_223 | (_ctrlsignals_T_225 | (_ctrlsignals_T_227 | (
    _ctrlsignals_T_229 | (_ctrlsignals_T_231 | _ctrlsignals_T_2296)))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2313 = _ctrlsignals_T_199 ? 1'h0 : _ctrlsignals_T_2312; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2314 = _ctrlsignals_T_197 ? 1'h0 : _ctrlsignals_T_2313; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2315 = _ctrlsignals_T_195 ? 1'h0 : _ctrlsignals_T_2314; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2316 = _ctrlsignals_T_193 ? 1'h0 : _ctrlsignals_T_2315; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2317 = _ctrlsignals_T_191 ? 1'h0 : _ctrlsignals_T_2316; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2318 = _ctrlsignals_T_189 ? 1'h0 : _ctrlsignals_T_2317; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2319 = _ctrlsignals_T_187 ? 1'h0 : _ctrlsignals_T_2318; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2320 = _ctrlsignals_T_185 ? 1'h0 : _ctrlsignals_T_2319; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2321 = _ctrlsignals_T_183 ? 1'h0 : _ctrlsignals_T_2320; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2322 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_2321; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2323 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_2322; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2324 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_2323; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2325 = _ctrlsignals_T_175 ? 1'h0 : _ctrlsignals_T_2324; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2326 = _ctrlsignals_T_173 ? 1'h0 : _ctrlsignals_T_2325; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2327 = _ctrlsignals_T_171 ? 1'h0 : _ctrlsignals_T_2326; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2328 = _ctrlsignals_T_169 ? 1'h0 : _ctrlsignals_T_2327; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2329 = _ctrlsignals_T_167 ? 1'h0 : _ctrlsignals_T_2328; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2330 = _ctrlsignals_T_165 ? 1'h0 : _ctrlsignals_T_2329; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2331 = _ctrlsignals_T_163 ? 1'h0 : _ctrlsignals_T_2330; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2332 = _ctrlsignals_T_161 ? 1'h0 : _ctrlsignals_T_2331; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2333 = _ctrlsignals_T_159 ? 1'h0 : _ctrlsignals_T_2332; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2334 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_2333; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2335 = _ctrlsignals_T_155 ? 1'h0 : _ctrlsignals_T_2334; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2336 = _ctrlsignals_T_153 ? 1'h0 : _ctrlsignals_T_2335; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2337 = _ctrlsignals_T_151 ? 1'h0 : _ctrlsignals_T_2336; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2338 = _ctrlsignals_T_149 ? 1'h0 : _ctrlsignals_T_2337; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2339 = _ctrlsignals_T_147 ? 1'h0 : _ctrlsignals_T_2338; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2340 = _ctrlsignals_T_145 ? 1'h0 : _ctrlsignals_T_2339; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2341 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_2340; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2342 = _ctrlsignals_T_141 ? 1'h0 : _ctrlsignals_T_2341; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2343 = _ctrlsignals_T_139 ? 1'h0 : _ctrlsignals_T_2342; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2344 = _ctrlsignals_T_137 ? 1'h0 : _ctrlsignals_T_2343; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2345 = _ctrlsignals_T_135 ? 1'h0 : _ctrlsignals_T_2344; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2346 = _ctrlsignals_T_133 ? 1'h0 : _ctrlsignals_T_2345; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2347 = _ctrlsignals_T_131 ? 1'h0 : _ctrlsignals_T_2346; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2348 = _ctrlsignals_T_129 ? 1'h0 : _ctrlsignals_T_2347; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2349 = _ctrlsignals_T_127 ? 1'h0 : _ctrlsignals_T_2348; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2350 = _ctrlsignals_T_125 ? 1'h0 : _ctrlsignals_T_2349; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2351 = _ctrlsignals_T_123 ? 1'h0 : _ctrlsignals_T_2350; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2352 = _ctrlsignals_T_121 ? 1'h0 : _ctrlsignals_T_2351; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2353 = _ctrlsignals_T_119 ? 1'h0 : _ctrlsignals_T_2352; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2354 = _ctrlsignals_T_117 ? 1'h0 : _ctrlsignals_T_2353; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2355 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_2354; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2356 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_2355; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2357 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_2356; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2358 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_2357; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2359 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_2358; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2360 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_2359; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2361 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_2360; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2362 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_2361; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2363 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_2362; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2364 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_2363; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2365 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_2364; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2366 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_2365; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2367 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_2366; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2368 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_2367; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2369 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_2368; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2370 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_2369; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2371 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_2370; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2372 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_2371; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2373 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_2372; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2374 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_2373; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2375 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_2374; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2376 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_2375; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2377 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_2376; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2378 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_2377; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2379 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_2378; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2380 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_2379; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2381 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_2380; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2382 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_2381; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2383 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_2382; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2384 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_2383; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2385 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_2384; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2386 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_2385; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2387 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_2386; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2388 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_2387; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2389 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_2388; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2390 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_2389; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2391 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_2390; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2392 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_2391; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2393 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_2392; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2394 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_2393; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2395 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_2394; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2396 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_2395; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2397 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_2396; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2398 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_2397; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2399 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_2398; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2400 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_2399; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2401 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_2400; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2402 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_2401; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2403 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_2402; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2404 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_2403; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2405 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_2404; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_2406 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_2405; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2563 = _ctrlsignals_T_181 ? 2'h3 : 2'h1; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2564 = _ctrlsignals_T_179 ? 2'h3 : _ctrlsignals_T_2563; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2565 = _ctrlsignals_T_177 ? 2'h3 : _ctrlsignals_T_2564; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2566 = _ctrlsignals_T_175 ? 2'h1 : _ctrlsignals_T_2565; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2567 = _ctrlsignals_T_173 ? 2'h1 : _ctrlsignals_T_2566; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2568 = _ctrlsignals_T_171 ? 2'h1 : _ctrlsignals_T_2567; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2569 = _ctrlsignals_T_169 ? 2'h1 : _ctrlsignals_T_2568; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2570 = _ctrlsignals_T_167 ? 2'h1 : _ctrlsignals_T_2569; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2571 = _ctrlsignals_T_165 ? 2'h1 : _ctrlsignals_T_2570; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2572 = _ctrlsignals_T_163 ? 2'h1 : _ctrlsignals_T_2571; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2573 = _ctrlsignals_T_161 ? 2'h1 : _ctrlsignals_T_2572; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2574 = _ctrlsignals_T_159 ? 2'h1 : _ctrlsignals_T_2573; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2575 = _ctrlsignals_T_143 ? 2'h1 : _ctrlsignals_T_2574; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2576 = _ctrlsignals_T_155 ? 2'h1 : _ctrlsignals_T_2575; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2577 = _ctrlsignals_T_153 ? 2'h1 : _ctrlsignals_T_2576; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2578 = _ctrlsignals_T_151 ? 2'h1 : _ctrlsignals_T_2577; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2579 = _ctrlsignals_T_149 ? 2'h1 : _ctrlsignals_T_2578; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2580 = _ctrlsignals_T_147 ? 2'h1 : _ctrlsignals_T_2579; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2581 = _ctrlsignals_T_145 ? 2'h1 : _ctrlsignals_T_2580; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2582 = _ctrlsignals_T_143 ? 2'h1 : _ctrlsignals_T_2581; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2583 = _ctrlsignals_T_141 ? 2'h1 : _ctrlsignals_T_2582; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2584 = _ctrlsignals_T_139 ? 2'h1 : _ctrlsignals_T_2583; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2585 = _ctrlsignals_T_137 ? 2'h1 : _ctrlsignals_T_2584; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2586 = _ctrlsignals_T_135 ? 2'h1 : _ctrlsignals_T_2585; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2587 = _ctrlsignals_T_133 ? 2'h1 : _ctrlsignals_T_2586; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2588 = _ctrlsignals_T_131 ? 2'h2 : _ctrlsignals_T_2587; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2589 = _ctrlsignals_T_129 ? 2'h2 : _ctrlsignals_T_2588; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2590 = _ctrlsignals_T_127 ? 2'h2 : _ctrlsignals_T_2589; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2591 = _ctrlsignals_T_125 ? 2'h2 : _ctrlsignals_T_2590; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2592 = _ctrlsignals_T_123 ? 2'h1 : _ctrlsignals_T_2591; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2593 = _ctrlsignals_T_121 ? 2'h1 : _ctrlsignals_T_2592; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2594 = _ctrlsignals_T_119 ? 2'h1 : _ctrlsignals_T_2593; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2595 = _ctrlsignals_T_117 ? 2'h1 : _ctrlsignals_T_2594; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2596 = _ctrlsignals_T_115 ? 2'h1 : _ctrlsignals_T_2595; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2597 = _ctrlsignals_T_113 ? 2'h1 : _ctrlsignals_T_2596; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2598 = _ctrlsignals_T_111 ? 2'h1 : _ctrlsignals_T_2597; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2599 = _ctrlsignals_T_109 ? 2'h1 : _ctrlsignals_T_2598; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2600 = _ctrlsignals_T_107 ? 2'h1 : _ctrlsignals_T_2599; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2601 = _ctrlsignals_T_105 ? 2'h1 : _ctrlsignals_T_2600; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2602 = _ctrlsignals_T_103 ? 2'h1 : _ctrlsignals_T_2601; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2603 = _ctrlsignals_T_101 ? 2'h1 : _ctrlsignals_T_2602; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2604 = _ctrlsignals_T_99 ? 2'h1 : _ctrlsignals_T_2603; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2605 = _ctrlsignals_T_97 ? 2'h1 : _ctrlsignals_T_2604; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2606 = _ctrlsignals_T_95 ? 2'h1 : _ctrlsignals_T_2605; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2607 = _ctrlsignals_T_93 ? 2'h1 : _ctrlsignals_T_2606; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2608 = _ctrlsignals_T_91 ? 2'h1 : _ctrlsignals_T_2607; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2609 = _ctrlsignals_T_89 ? 2'h1 : _ctrlsignals_T_2608; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2610 = _ctrlsignals_T_87 ? 2'h1 : _ctrlsignals_T_2609; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2611 = _ctrlsignals_T_85 ? 2'h1 : _ctrlsignals_T_2610; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2612 = _ctrlsignals_T_83 ? 2'h1 : _ctrlsignals_T_2611; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2613 = _ctrlsignals_T_81 ? 2'h1 : _ctrlsignals_T_2612; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2614 = _ctrlsignals_T_79 ? 2'h1 : _ctrlsignals_T_2613; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2615 = _ctrlsignals_T_77 ? 2'h1 : _ctrlsignals_T_2614; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2616 = _ctrlsignals_T_75 ? 2'h1 : _ctrlsignals_T_2615; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2617 = _ctrlsignals_T_73 ? 2'h1 : _ctrlsignals_T_2616; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2618 = _ctrlsignals_T_71 ? 2'h1 : _ctrlsignals_T_2617; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2619 = _ctrlsignals_T_69 ? 2'h1 : _ctrlsignals_T_2618; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2620 = _ctrlsignals_T_67 ? 2'h1 : _ctrlsignals_T_2619; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2621 = _ctrlsignals_T_65 ? 2'h3 : _ctrlsignals_T_2620; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2622 = _ctrlsignals_T_63 ? 2'h3 : _ctrlsignals_T_2621; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2623 = _ctrlsignals_T_61 ? 2'h3 : _ctrlsignals_T_2622; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2624 = _ctrlsignals_T_59 ? 2'h1 : _ctrlsignals_T_2623; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2625 = _ctrlsignals_T_57 ? 2'h1 : _ctrlsignals_T_2624; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2626 = _ctrlsignals_T_55 ? 2'h1 : _ctrlsignals_T_2625; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2627 = _ctrlsignals_T_53 ? 2'h1 : _ctrlsignals_T_2626; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2628 = _ctrlsignals_T_51 ? 2'h1 : _ctrlsignals_T_2627; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2629 = _ctrlsignals_T_49 ? 2'h1 : _ctrlsignals_T_2628; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2630 = _ctrlsignals_T_47 ? 2'h1 : _ctrlsignals_T_2629; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2631 = _ctrlsignals_T_45 ? 2'h1 : _ctrlsignals_T_2630; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2632 = _ctrlsignals_T_43 ? 2'h1 : _ctrlsignals_T_2631; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2633 = _ctrlsignals_T_41 ? 2'h1 : _ctrlsignals_T_2632; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2634 = _ctrlsignals_T_39 ? 2'h1 : _ctrlsignals_T_2633; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2635 = _ctrlsignals_T_37 ? 2'h1 : _ctrlsignals_T_2634; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2636 = _ctrlsignals_T_35 ? 2'h1 : _ctrlsignals_T_2635; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2637 = _ctrlsignals_T_33 ? 2'h0 : _ctrlsignals_T_2636; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2638 = _ctrlsignals_T_31 ? 2'h0 : _ctrlsignals_T_2637; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2639 = _ctrlsignals_T_29 ? 2'h0 : _ctrlsignals_T_2638; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2640 = _ctrlsignals_T_27 ? 2'h0 : _ctrlsignals_T_2639; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2641 = _ctrlsignals_T_25 ? 2'h0 : _ctrlsignals_T_2640; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2642 = _ctrlsignals_T_23 ? 2'h0 : _ctrlsignals_T_2641; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2643 = _ctrlsignals_T_21 ? 2'h0 : _ctrlsignals_T_2642; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2644 = _ctrlsignals_T_19 ? 2'h0 : _ctrlsignals_T_2643; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2645 = _ctrlsignals_T_17 ? 2'h1 : _ctrlsignals_T_2644; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2646 = _ctrlsignals_T_15 ? 2'h1 : _ctrlsignals_T_2645; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2647 = _ctrlsignals_T_13 ? 2'h0 : _ctrlsignals_T_2646; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2648 = _ctrlsignals_T_11 ? 2'h0 : _ctrlsignals_T_2647; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2649 = _ctrlsignals_T_9 ? 2'h0 : _ctrlsignals_T_2648; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2650 = _ctrlsignals_T_7 ? 2'h0 : _ctrlsignals_T_2649; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2651 = _ctrlsignals_T_5 ? 2'h0 : _ctrlsignals_T_2650; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2652 = _ctrlsignals_T_3 ? 2'h0 : _ctrlsignals_T_2651; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2656 = _ctrlsignals_T_477 ? 2'h2 : 2'h1; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2657 = _ctrlsignals_T_475 ? 2'h1 : _ctrlsignals_T_2656; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2658 = _ctrlsignals_T_473 ? 2'h1 : _ctrlsignals_T_2657; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2659 = _ctrlsignals_T_471 ? 2'h1 : _ctrlsignals_T_2658; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2660 = _ctrlsignals_T_469 ? 2'h1 : _ctrlsignals_T_2659; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2661 = _ctrlsignals_T_467 ? 2'h2 : _ctrlsignals_T_2660; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2662 = _ctrlsignals_T_465 ? 2'h2 : _ctrlsignals_T_2661; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2663 = _ctrlsignals_T_463 ? 2'h2 : _ctrlsignals_T_2662; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2664 = _ctrlsignals_T_461 ? 2'h2 : _ctrlsignals_T_2663; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2665 = _ctrlsignals_T_459 ? 2'h2 : _ctrlsignals_T_2664; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2666 = _ctrlsignals_T_445 ? 2'h2 : _ctrlsignals_T_2665; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2667 = _ctrlsignals_T_443 ? 2'h2 : _ctrlsignals_T_2666; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2668 = _ctrlsignals_T_453 ? 2'h2 : _ctrlsignals_T_2667; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2669 = _ctrlsignals_T_451 ? 2'h2 : _ctrlsignals_T_2668; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2670 = _ctrlsignals_T_449 ? 2'h2 : _ctrlsignals_T_2669; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2671 = _ctrlsignals_T_447 ? 2'h2 : _ctrlsignals_T_2670; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2672 = _ctrlsignals_T_445 ? 2'h2 : _ctrlsignals_T_2671; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2673 = _ctrlsignals_T_443 ? 2'h2 : _ctrlsignals_T_2672; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2674 = _ctrlsignals_T_441 ? 2'h2 : _ctrlsignals_T_2673; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2675 = _ctrlsignals_T_439 ? 2'h2 : _ctrlsignals_T_2674; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2676 = _ctrlsignals_T_437 ? 2'h2 : _ctrlsignals_T_2675; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2677 = _ctrlsignals_T_435 ? 2'h2 : _ctrlsignals_T_2676; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2678 = _ctrlsignals_T_433 ? 2'h2 : _ctrlsignals_T_2677; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2679 = _ctrlsignals_T_431 ? 2'h2 : _ctrlsignals_T_2678; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2680 = _ctrlsignals_T_429 ? 2'h2 : _ctrlsignals_T_2679; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2681 = _ctrlsignals_T_427 ? 2'h2 : _ctrlsignals_T_2680; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2682 = _ctrlsignals_T_425 ? 2'h2 : _ctrlsignals_T_2681; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2683 = _ctrlsignals_T_423 ? 2'h2 : _ctrlsignals_T_2682; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2684 = _ctrlsignals_T_421 ? 2'h2 : _ctrlsignals_T_2683; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2685 = _ctrlsignals_T_419 ? 2'h2 : _ctrlsignals_T_2684; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2686 = _ctrlsignals_T_417 ? 2'h2 : _ctrlsignals_T_2685; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2687 = _ctrlsignals_T_415 ? 2'h2 : _ctrlsignals_T_2686; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2688 = _ctrlsignals_T_413 ? 2'h2 : _ctrlsignals_T_2687; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2689 = _ctrlsignals_T_411 ? 2'h2 : _ctrlsignals_T_2688; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2690 = _ctrlsignals_T_409 ? 2'h2 : _ctrlsignals_T_2689; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2691 = _ctrlsignals_T_407 ? 2'h2 : _ctrlsignals_T_2690; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2692 = _ctrlsignals_T_405 ? 2'h2 : _ctrlsignals_T_2691; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2693 = _ctrlsignals_T_403 ? 2'h2 : _ctrlsignals_T_2692; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2694 = _ctrlsignals_T_401 ? 2'h2 : _ctrlsignals_T_2693; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2695 = _ctrlsignals_T_399 ? 2'h2 : _ctrlsignals_T_2694; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2696 = _ctrlsignals_T_397 ? 2'h2 : _ctrlsignals_T_2695; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2697 = _ctrlsignals_T_395 ? 2'h2 : _ctrlsignals_T_2696; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2698 = _ctrlsignals_T_393 ? 2'h2 : _ctrlsignals_T_2697; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2699 = _ctrlsignals_T_391 ? 2'h2 : _ctrlsignals_T_2698; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2700 = _ctrlsignals_T_389 ? 2'h2 : _ctrlsignals_T_2699; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2701 = _ctrlsignals_T_387 ? 2'h2 : _ctrlsignals_T_2700; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2702 = _ctrlsignals_T_385 ? 2'h2 : _ctrlsignals_T_2701; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2703 = _ctrlsignals_T_383 ? 2'h2 : _ctrlsignals_T_2702; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2704 = _ctrlsignals_T_381 ? 2'h2 : _ctrlsignals_T_2703; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2705 = _ctrlsignals_T_379 ? 2'h2 : _ctrlsignals_T_2704; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2706 = _ctrlsignals_T_377 ? 2'h2 : _ctrlsignals_T_2705; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2707 = _ctrlsignals_T_375 ? 2'h2 : _ctrlsignals_T_2706; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2708 = _ctrlsignals_T_373 ? 2'h2 : _ctrlsignals_T_2707; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2709 = _ctrlsignals_T_371 ? 2'h2 : _ctrlsignals_T_2708; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2710 = _ctrlsignals_T_369 ? 2'h2 : _ctrlsignals_T_2709; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2711 = _ctrlsignals_T_367 ? 2'h2 : _ctrlsignals_T_2710; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2712 = _ctrlsignals_T_365 ? 2'h2 : _ctrlsignals_T_2711; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2713 = _ctrlsignals_T_363 ? 2'h1 : _ctrlsignals_T_2712; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2714 = _ctrlsignals_T_361 ? 2'h2 : _ctrlsignals_T_2713; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2715 = _ctrlsignals_T_359 ? 2'h2 : _ctrlsignals_T_2714; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2716 = _ctrlsignals_T_357 ? 2'h2 : _ctrlsignals_T_2715; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2717 = _ctrlsignals_T_355 ? 2'h2 : _ctrlsignals_T_2716; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2718 = _ctrlsignals_T_353 ? 2'h2 : _ctrlsignals_T_2717; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2719 = _ctrlsignals_T_351 ? 2'h2 : _ctrlsignals_T_2718; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2720 = _ctrlsignals_T_349 ? 2'h2 : _ctrlsignals_T_2719; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2721 = _ctrlsignals_T_347 ? 2'h2 : _ctrlsignals_T_2720; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2722 = _ctrlsignals_T_345 ? 2'h2 : _ctrlsignals_T_2721; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2723 = _ctrlsignals_T_343 ? 2'h2 : _ctrlsignals_T_2722; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2724 = _ctrlsignals_T_341 ? 2'h2 : _ctrlsignals_T_2723; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2725 = _ctrlsignals_T_339 ? 2'h2 : _ctrlsignals_T_2724; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2726 = _ctrlsignals_T_337 ? 2'h2 : _ctrlsignals_T_2725; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2727 = _ctrlsignals_T_335 ? 2'h2 : _ctrlsignals_T_2726; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2728 = _ctrlsignals_T_333 ? 2'h2 : _ctrlsignals_T_2727; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2729 = _ctrlsignals_T_331 ? 2'h2 : _ctrlsignals_T_2728; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2730 = _ctrlsignals_T_329 ? 2'h2 : _ctrlsignals_T_2729; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2731 = _ctrlsignals_T_327 ? 2'h2 : _ctrlsignals_T_2730; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2732 = _ctrlsignals_T_325 ? 2'h2 : _ctrlsignals_T_2731; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2733 = _ctrlsignals_T_323 ? 2'h2 : _ctrlsignals_T_2732; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2734 = _ctrlsignals_T_321 ? 2'h2 : _ctrlsignals_T_2733; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2735 = _ctrlsignals_T_319 ? 2'h2 : _ctrlsignals_T_2734; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2736 = _ctrlsignals_T_317 ? 2'h2 : _ctrlsignals_T_2735; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2737 = _ctrlsignals_T_315 ? 2'h2 : _ctrlsignals_T_2736; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2738 = _ctrlsignals_T_313 ? 2'h2 : _ctrlsignals_T_2737; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2739 = _ctrlsignals_T_311 ? 2'h2 : _ctrlsignals_T_2738; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2740 = _ctrlsignals_T_309 ? 2'h2 : _ctrlsignals_T_2739; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2741 = _ctrlsignals_T_307 ? 2'h2 : _ctrlsignals_T_2740; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2742 = _ctrlsignals_T_305 ? 2'h2 : _ctrlsignals_T_2741; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2743 = _ctrlsignals_T_303 ? 2'h2 : _ctrlsignals_T_2742; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2744 = _ctrlsignals_T_301 ? 2'h2 : _ctrlsignals_T_2743; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2745 = _ctrlsignals_T_299 ? 2'h2 : _ctrlsignals_T_2744; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2746 = _ctrlsignals_T_297 ? 2'h2 : _ctrlsignals_T_2745; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2747 = _ctrlsignals_T_295 ? 2'h2 : _ctrlsignals_T_2746; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2748 = _ctrlsignals_T_293 ? 2'h2 : _ctrlsignals_T_2747; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2749 = _ctrlsignals_T_291 ? 2'h2 : _ctrlsignals_T_2748; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2750 = _ctrlsignals_T_289 ? 2'h2 : _ctrlsignals_T_2749; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2751 = _ctrlsignals_T_287 ? 2'h2 : _ctrlsignals_T_2750; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2752 = _ctrlsignals_T_285 ? 2'h2 : _ctrlsignals_T_2751; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2753 = _ctrlsignals_T_283 ? 2'h2 : _ctrlsignals_T_2752; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2754 = _ctrlsignals_T_281 ? 2'h2 : _ctrlsignals_T_2753; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2755 = _ctrlsignals_T_279 ? 2'h2 : _ctrlsignals_T_2754; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2756 = _ctrlsignals_T_277 ? 2'h2 : _ctrlsignals_T_2755; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2757 = _ctrlsignals_T_275 ? 2'h2 : _ctrlsignals_T_2756; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2758 = _ctrlsignals_T_273 ? 2'h2 : _ctrlsignals_T_2757; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2759 = _ctrlsignals_T_271 ? 2'h2 : _ctrlsignals_T_2758; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2760 = _ctrlsignals_T_269 ? 2'h2 : _ctrlsignals_T_2759; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2761 = _ctrlsignals_T_267 ? 2'h2 : _ctrlsignals_T_2760; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2762 = _ctrlsignals_T_265 ? 2'h2 : _ctrlsignals_T_2761; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2763 = _ctrlsignals_T_263 ? 2'h2 : _ctrlsignals_T_2762; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2764 = _ctrlsignals_T_261 ? 2'h2 : _ctrlsignals_T_2763; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2765 = _ctrlsignals_T_259 ? 2'h2 : _ctrlsignals_T_2764; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2766 = _ctrlsignals_T_257 ? 2'h2 : _ctrlsignals_T_2765; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2767 = _ctrlsignals_T_255 ? 2'h2 : _ctrlsignals_T_2766; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2768 = _ctrlsignals_T_253 ? 2'h2 : _ctrlsignals_T_2767; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2769 = _ctrlsignals_T_251 ? 2'h2 : _ctrlsignals_T_2768; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2770 = _ctrlsignals_T_249 ? 2'h2 : _ctrlsignals_T_2769; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2771 = _ctrlsignals_T_247 ? 2'h2 : _ctrlsignals_T_2770; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2772 = _ctrlsignals_T_245 ? 2'h2 : _ctrlsignals_T_2771; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2773 = _ctrlsignals_T_243 ? 2'h2 : _ctrlsignals_T_2772; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2774 = _ctrlsignals_T_241 ? 2'h2 : _ctrlsignals_T_2773; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2775 = _ctrlsignals_T_239 ? 2'h2 : _ctrlsignals_T_2774; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2776 = _ctrlsignals_T_237 ? 2'h2 : _ctrlsignals_T_2775; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2777 = _ctrlsignals_T_235 ? 2'h2 : _ctrlsignals_T_2776; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2778 = _ctrlsignals_T_233 ? 2'h2 : _ctrlsignals_T_2777; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2779 = _ctrlsignals_T_231 ? 2'h2 : _ctrlsignals_T_2778; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2780 = _ctrlsignals_T_229 ? 2'h2 : _ctrlsignals_T_2779; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2781 = _ctrlsignals_T_227 ? 2'h2 : _ctrlsignals_T_2780; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2782 = _ctrlsignals_T_225 ? 2'h2 : _ctrlsignals_T_2781; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2783 = _ctrlsignals_T_223 ? 2'h2 : _ctrlsignals_T_2782; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2784 = _ctrlsignals_T_221 ? 2'h2 : _ctrlsignals_T_2783; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2785 = _ctrlsignals_T_219 ? 2'h2 : _ctrlsignals_T_2784; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2786 = _ctrlsignals_T_217 ? 2'h2 : _ctrlsignals_T_2785; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2787 = _ctrlsignals_T_215 ? 2'h2 : _ctrlsignals_T_2786; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2788 = _ctrlsignals_T_213 ? 2'h2 : _ctrlsignals_T_2787; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2789 = _ctrlsignals_T_211 ? 2'h2 : _ctrlsignals_T_2788; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2790 = _ctrlsignals_T_209 ? 2'h2 : _ctrlsignals_T_2789; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2791 = _ctrlsignals_T_207 ? 2'h2 : _ctrlsignals_T_2790; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2792 = _ctrlsignals_T_205 ? 2'h2 : _ctrlsignals_T_2791; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2793 = _ctrlsignals_T_203 ? 2'h2 : _ctrlsignals_T_2792; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2794 = _ctrlsignals_T_201 ? 2'h2 : _ctrlsignals_T_2793; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2795 = _ctrlsignals_T_199 ? 2'h2 : _ctrlsignals_T_2794; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2796 = _ctrlsignals_T_197 ? 2'h2 : _ctrlsignals_T_2795; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2797 = _ctrlsignals_T_195 ? 2'h2 : _ctrlsignals_T_2796; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2798 = _ctrlsignals_T_193 ? 2'h2 : _ctrlsignals_T_2797; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2799 = _ctrlsignals_T_191 ? 2'h2 : _ctrlsignals_T_2798; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2800 = _ctrlsignals_T_189 ? 2'h2 : _ctrlsignals_T_2799; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2801 = _ctrlsignals_T_187 ? 2'h2 : _ctrlsignals_T_2800; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2802 = _ctrlsignals_T_185 ? 2'h2 : _ctrlsignals_T_2801; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2803 = _ctrlsignals_T_183 ? 2'h2 : _ctrlsignals_T_2802; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2804 = _ctrlsignals_T_181 ? 2'h2 : _ctrlsignals_T_2803; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2805 = _ctrlsignals_T_179 ? 2'h1 : _ctrlsignals_T_2804; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2806 = _ctrlsignals_T_177 ? 2'h1 : _ctrlsignals_T_2805; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2807 = _ctrlsignals_T_175 ? 2'h2 : _ctrlsignals_T_2806; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2808 = _ctrlsignals_T_173 ? 2'h1 : _ctrlsignals_T_2807; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2809 = _ctrlsignals_T_171 ? 2'h1 : _ctrlsignals_T_2808; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2810 = _ctrlsignals_T_169 ? 2'h1 : _ctrlsignals_T_2809; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2811 = _ctrlsignals_T_167 ? 2'h1 : _ctrlsignals_T_2810; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2812 = _ctrlsignals_T_165 ? 2'h1 : _ctrlsignals_T_2811; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2813 = _ctrlsignals_T_163 ? 2'h1 : _ctrlsignals_T_2812; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2814 = _ctrlsignals_T_161 ? 2'h1 : _ctrlsignals_T_2813; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2815 = _ctrlsignals_T_159 ? 2'h1 : _ctrlsignals_T_2814; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2816 = _ctrlsignals_T_143 ? 2'h1 : _ctrlsignals_T_2815; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2817 = _ctrlsignals_T_155 ? 2'h1 : _ctrlsignals_T_2816; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2818 = _ctrlsignals_T_153 ? 2'h1 : _ctrlsignals_T_2817; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2819 = _ctrlsignals_T_151 ? 2'h1 : _ctrlsignals_T_2818; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2820 = _ctrlsignals_T_149 ? 2'h1 : _ctrlsignals_T_2819; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2821 = _ctrlsignals_T_147 ? 2'h1 : _ctrlsignals_T_2820; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2822 = _ctrlsignals_T_145 ? 2'h1 : _ctrlsignals_T_2821; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2823 = _ctrlsignals_T_143 ? 2'h1 : _ctrlsignals_T_2822; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2824 = _ctrlsignals_T_141 ? 2'h1 : _ctrlsignals_T_2823; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2825 = _ctrlsignals_T_139 ? 2'h1 : _ctrlsignals_T_2824; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2826 = _ctrlsignals_T_137 ? 2'h1 : _ctrlsignals_T_2825; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2827 = _ctrlsignals_T_135 ? 2'h1 : _ctrlsignals_T_2826; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2828 = _ctrlsignals_T_133 ? 2'h1 : _ctrlsignals_T_2827; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2829 = _ctrlsignals_T_131 ? 2'h1 : _ctrlsignals_T_2828; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2830 = _ctrlsignals_T_129 ? 2'h1 : _ctrlsignals_T_2829; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2831 = _ctrlsignals_T_127 ? 2'h1 : _ctrlsignals_T_2830; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2832 = _ctrlsignals_T_125 ? 2'h1 : _ctrlsignals_T_2831; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2833 = _ctrlsignals_T_123 ? 2'h1 : _ctrlsignals_T_2832; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2834 = _ctrlsignals_T_121 ? 2'h1 : _ctrlsignals_T_2833; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2835 = _ctrlsignals_T_119 ? 2'h1 : _ctrlsignals_T_2834; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2836 = _ctrlsignals_T_117 ? 2'h1 : _ctrlsignals_T_2835; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2837 = _ctrlsignals_T_115 ? 2'h1 : _ctrlsignals_T_2836; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2838 = _ctrlsignals_T_113 ? 2'h1 : _ctrlsignals_T_2837; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2839 = _ctrlsignals_T_111 ? 2'h1 : _ctrlsignals_T_2838; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2840 = _ctrlsignals_T_109 ? 2'h1 : _ctrlsignals_T_2839; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2841 = _ctrlsignals_T_107 ? 2'h3 : _ctrlsignals_T_2840; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2842 = _ctrlsignals_T_105 ? 2'h3 : _ctrlsignals_T_2841; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2843 = _ctrlsignals_T_103 ? 2'h3 : _ctrlsignals_T_2842; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2844 = _ctrlsignals_T_101 ? 2'h3 : _ctrlsignals_T_2843; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2845 = _ctrlsignals_T_99 ? 2'h1 : _ctrlsignals_T_2844; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2846 = _ctrlsignals_T_97 ? 2'h1 : _ctrlsignals_T_2845; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2847 = _ctrlsignals_T_95 ? 2'h1 : _ctrlsignals_T_2846; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2848 = _ctrlsignals_T_93 ? 2'h1 : _ctrlsignals_T_2847; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2849 = _ctrlsignals_T_91 ? 2'h1 : _ctrlsignals_T_2848; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2850 = _ctrlsignals_T_89 ? 2'h1 : _ctrlsignals_T_2849; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2851 = _ctrlsignals_T_87 ? 2'h1 : _ctrlsignals_T_2850; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2852 = _ctrlsignals_T_85 ? 2'h1 : _ctrlsignals_T_2851; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2853 = _ctrlsignals_T_83 ? 2'h1 : _ctrlsignals_T_2852; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2854 = _ctrlsignals_T_81 ? 2'h1 : _ctrlsignals_T_2853; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2855 = _ctrlsignals_T_79 ? 2'h3 : _ctrlsignals_T_2854; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2856 = _ctrlsignals_T_77 ? 2'h3 : _ctrlsignals_T_2855; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2857 = _ctrlsignals_T_75 ? 2'h3 : _ctrlsignals_T_2856; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2858 = _ctrlsignals_T_73 ? 2'h3 : _ctrlsignals_T_2857; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2859 = _ctrlsignals_T_71 ? 2'h3 : _ctrlsignals_T_2858; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2860 = _ctrlsignals_T_69 ? 2'h3 : _ctrlsignals_T_2859; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2861 = _ctrlsignals_T_67 ? 2'h3 : _ctrlsignals_T_2860; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2862 = _ctrlsignals_T_65 ? 2'h3 : _ctrlsignals_T_2861; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2863 = _ctrlsignals_T_63 ? 2'h3 : _ctrlsignals_T_2862; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2864 = _ctrlsignals_T_61 ? 2'h3 : _ctrlsignals_T_2863; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2865 = _ctrlsignals_T_59 ? 2'h3 : _ctrlsignals_T_2864; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2866 = _ctrlsignals_T_57 ? 2'h3 : _ctrlsignals_T_2865; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2867 = _ctrlsignals_T_55 ? 2'h3 : _ctrlsignals_T_2866; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2868 = _ctrlsignals_T_53 ? 2'h3 : _ctrlsignals_T_2867; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2869 = _ctrlsignals_T_51 ? 2'h3 : _ctrlsignals_T_2868; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2870 = _ctrlsignals_T_49 ? 2'h1 : _ctrlsignals_T_2869; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2871 = _ctrlsignals_T_47 ? 2'h1 : _ctrlsignals_T_2870; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2872 = _ctrlsignals_T_45 ? 2'h1 : _ctrlsignals_T_2871; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2873 = _ctrlsignals_T_43 ? 2'h1 : _ctrlsignals_T_2872; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2874 = _ctrlsignals_T_41 ? 2'h1 : _ctrlsignals_T_2873; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2875 = _ctrlsignals_T_39 ? 2'h1 : _ctrlsignals_T_2874; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2876 = _ctrlsignals_T_37 ? 2'h1 : _ctrlsignals_T_2875; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2877 = _ctrlsignals_T_35 ? 2'h3 : _ctrlsignals_T_2876; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2878 = _ctrlsignals_T_33 ? 2'h0 : _ctrlsignals_T_2877; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2879 = _ctrlsignals_T_31 ? 2'h0 : _ctrlsignals_T_2878; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2880 = _ctrlsignals_T_29 ? 2'h1 : _ctrlsignals_T_2879; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2881 = _ctrlsignals_T_27 ? 2'h1 : _ctrlsignals_T_2880; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2882 = _ctrlsignals_T_25 ? 2'h1 : _ctrlsignals_T_2881; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2883 = _ctrlsignals_T_23 ? 2'h1 : _ctrlsignals_T_2882; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2884 = _ctrlsignals_T_21 ? 2'h1 : _ctrlsignals_T_2883; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2885 = _ctrlsignals_T_19 ? 2'h1 : _ctrlsignals_T_2884; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2886 = _ctrlsignals_T_17 ? 2'h1 : _ctrlsignals_T_2885; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2887 = _ctrlsignals_T_15 ? 2'h2 : _ctrlsignals_T_2886; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2888 = _ctrlsignals_T_13 ? 2'h1 : _ctrlsignals_T_2887; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2889 = _ctrlsignals_T_11 ? 2'h2 : _ctrlsignals_T_2888; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2890 = _ctrlsignals_T_9 ? 2'h2 : _ctrlsignals_T_2889; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2891 = _ctrlsignals_T_7 ? 2'h2 : _ctrlsignals_T_2890; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2892 = _ctrlsignals_T_5 ? 2'h2 : _ctrlsignals_T_2891; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2893 = _ctrlsignals_T_3 ? 2'h2 : _ctrlsignals_T_2892; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2895 = _ctrlsignals_T_481 ? 2'h3 : 2'h1; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2896 = _ctrlsignals_T_479 ? 2'h1 : _ctrlsignals_T_2895; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2897 = _ctrlsignals_T_477 ? 2'h1 : _ctrlsignals_T_2896; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2898 = _ctrlsignals_T_475 ? 2'h1 : _ctrlsignals_T_2897; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2899 = _ctrlsignals_T_473 ? 2'h3 : _ctrlsignals_T_2898; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2900 = _ctrlsignals_T_471 ? 2'h1 : _ctrlsignals_T_2899; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2901 = _ctrlsignals_T_469 ? 2'h2 : _ctrlsignals_T_2900; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2902 = _ctrlsignals_T_467 ? 2'h1 : _ctrlsignals_T_2901; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2903 = _ctrlsignals_T_465 ? 2'h1 : _ctrlsignals_T_2902; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2904 = _ctrlsignals_T_463 ? 2'h1 : _ctrlsignals_T_2903; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2905 = _ctrlsignals_T_461 ? 2'h1 : _ctrlsignals_T_2904; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2906 = _ctrlsignals_T_459 ? 2'h1 : _ctrlsignals_T_2905; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2907 = _ctrlsignals_T_445 ? 2'h1 : _ctrlsignals_T_2906; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2908 = _ctrlsignals_T_443 ? 2'h2 : _ctrlsignals_T_2907; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2909 = _ctrlsignals_T_453 ? 2'h1 : _ctrlsignals_T_2908; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2910 = _ctrlsignals_T_451 ? 2'h2 : _ctrlsignals_T_2909; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2911 = _ctrlsignals_T_449 ? 2'h1 : _ctrlsignals_T_2910; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2912 = _ctrlsignals_T_447 ? 2'h2 : _ctrlsignals_T_2911; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2913 = _ctrlsignals_T_445 ? 2'h1 : _ctrlsignals_T_2912; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2914 = _ctrlsignals_T_443 ? 2'h2 : _ctrlsignals_T_2913; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2915 = _ctrlsignals_T_441 ? 2'h1 : _ctrlsignals_T_2914; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2916 = _ctrlsignals_T_439 ? 2'h1 : _ctrlsignals_T_2915; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2917 = _ctrlsignals_T_437 ? 2'h1 : _ctrlsignals_T_2916; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2918 = _ctrlsignals_T_435 ? 2'h1 : _ctrlsignals_T_2917; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2919 = _ctrlsignals_T_433 ? 2'h2 : _ctrlsignals_T_2918; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2920 = _ctrlsignals_T_431 ? 2'h2 : _ctrlsignals_T_2919; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2921 = _ctrlsignals_T_429 ? 2'h2 : _ctrlsignals_T_2920; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2922 = _ctrlsignals_T_427 ? 2'h2 : _ctrlsignals_T_2921; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2923 = _ctrlsignals_T_425 ? 2'h1 : _ctrlsignals_T_2922; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2924 = _ctrlsignals_T_423 ? 2'h1 : _ctrlsignals_T_2923; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2925 = _ctrlsignals_T_421 ? 2'h1 : _ctrlsignals_T_2924; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2926 = _ctrlsignals_T_419 ? 2'h2 : _ctrlsignals_T_2925; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2927 = _ctrlsignals_T_417 ? 2'h1 : _ctrlsignals_T_2926; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2928 = _ctrlsignals_T_415 ? 2'h2 : _ctrlsignals_T_2927; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2929 = _ctrlsignals_T_413 ? 2'h1 : _ctrlsignals_T_2928; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2930 = _ctrlsignals_T_411 ? 2'h2 : _ctrlsignals_T_2929; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2931 = _ctrlsignals_T_409 ? 2'h1 : _ctrlsignals_T_2930; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2932 = _ctrlsignals_T_407 ? 2'h2 : _ctrlsignals_T_2931; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2933 = _ctrlsignals_T_405 ? 2'h1 : _ctrlsignals_T_2932; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2934 = _ctrlsignals_T_403 ? 2'h2 : _ctrlsignals_T_2933; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2935 = _ctrlsignals_T_401 ? 2'h1 : _ctrlsignals_T_2934; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2936 = _ctrlsignals_T_399 ? 2'h2 : _ctrlsignals_T_2935; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2937 = _ctrlsignals_T_397 ? 2'h1 : _ctrlsignals_T_2936; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2938 = _ctrlsignals_T_395 ? 2'h2 : _ctrlsignals_T_2937; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2939 = _ctrlsignals_T_393 ? 2'h1 : _ctrlsignals_T_2938; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2940 = _ctrlsignals_T_391 ? 2'h2 : _ctrlsignals_T_2939; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2941 = _ctrlsignals_T_389 ? 2'h1 : _ctrlsignals_T_2940; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2942 = _ctrlsignals_T_387 ? 2'h2 : _ctrlsignals_T_2941; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2943 = _ctrlsignals_T_385 ? 2'h1 : _ctrlsignals_T_2942; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2944 = _ctrlsignals_T_383 ? 2'h2 : _ctrlsignals_T_2943; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2945 = _ctrlsignals_T_381 ? 2'h1 : _ctrlsignals_T_2944; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2946 = _ctrlsignals_T_379 ? 2'h2 : _ctrlsignals_T_2945; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2947 = _ctrlsignals_T_377 ? 2'h1 : _ctrlsignals_T_2946; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2948 = _ctrlsignals_T_375 ? 2'h2 : _ctrlsignals_T_2947; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2949 = _ctrlsignals_T_373 ? 2'h1 : _ctrlsignals_T_2948; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2950 = _ctrlsignals_T_371 ? 2'h2 : _ctrlsignals_T_2949; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2951 = _ctrlsignals_T_369 ? 2'h3 : _ctrlsignals_T_2950; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2952 = _ctrlsignals_T_367 ? 2'h1 : _ctrlsignals_T_2951; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2953 = _ctrlsignals_T_365 ? 2'h2 : _ctrlsignals_T_2952; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2954 = _ctrlsignals_T_363 ? 2'h1 : _ctrlsignals_T_2953; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2955 = _ctrlsignals_T_361 ? 2'h2 : _ctrlsignals_T_2954; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2956 = _ctrlsignals_T_359 ? 2'h2 : _ctrlsignals_T_2955; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2957 = _ctrlsignals_T_357 ? 2'h2 : _ctrlsignals_T_2956; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2958 = _ctrlsignals_T_355 ? 2'h2 : _ctrlsignals_T_2957; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2959 = _ctrlsignals_T_353 ? 2'h2 : _ctrlsignals_T_2958; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2960 = _ctrlsignals_T_351 ? 2'h2 : _ctrlsignals_T_2959; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2961 = _ctrlsignals_T_349 ? 2'h2 : _ctrlsignals_T_2960; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2962 = _ctrlsignals_T_347 ? 2'h2 : _ctrlsignals_T_2961; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2963 = _ctrlsignals_T_345 ? 2'h2 : _ctrlsignals_T_2962; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2964 = _ctrlsignals_T_343 ? 2'h3 : _ctrlsignals_T_2963; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2965 = _ctrlsignals_T_341 ? 2'h2 : _ctrlsignals_T_2964; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2966 = _ctrlsignals_T_339 ? 2'h3 : _ctrlsignals_T_2965; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2967 = _ctrlsignals_T_337 ? 2'h1 : _ctrlsignals_T_2966; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2968 = _ctrlsignals_T_335 ? 2'h3 : _ctrlsignals_T_2967; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2969 = _ctrlsignals_T_333 ? 2'h2 : _ctrlsignals_T_2968; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2970 = _ctrlsignals_T_331 ? 2'h1 : _ctrlsignals_T_2969; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2971 = _ctrlsignals_T_329 ? 2'h3 : _ctrlsignals_T_2970; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2972 = _ctrlsignals_T_327 ? 2'h2 : _ctrlsignals_T_2971; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2973 = _ctrlsignals_T_325 ? 2'h3 : _ctrlsignals_T_2972; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2974 = _ctrlsignals_T_323 ? 2'h1 : _ctrlsignals_T_2973; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2975 = _ctrlsignals_T_321 ? 2'h2 : _ctrlsignals_T_2974; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2976 = _ctrlsignals_T_319 ? 2'h3 : _ctrlsignals_T_2975; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2977 = _ctrlsignals_T_317 ? 2'h1 : _ctrlsignals_T_2976; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2978 = _ctrlsignals_T_315 ? 2'h2 : _ctrlsignals_T_2977; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2979 = _ctrlsignals_T_313 ? 2'h3 : _ctrlsignals_T_2978; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2980 = _ctrlsignals_T_311 ? 2'h1 : _ctrlsignals_T_2979; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2981 = _ctrlsignals_T_309 ? 2'h2 : _ctrlsignals_T_2980; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2982 = _ctrlsignals_T_307 ? 2'h1 : _ctrlsignals_T_2981; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2983 = _ctrlsignals_T_305 ? 2'h1 : _ctrlsignals_T_2982; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2984 = _ctrlsignals_T_303 ? 2'h1 : _ctrlsignals_T_2983; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2985 = _ctrlsignals_T_301 ? 2'h2 : _ctrlsignals_T_2984; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2986 = _ctrlsignals_T_299 ? 2'h1 : _ctrlsignals_T_2985; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2987 = _ctrlsignals_T_297 ? 2'h2 : _ctrlsignals_T_2986; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2988 = _ctrlsignals_T_295 ? 2'h1 : _ctrlsignals_T_2987; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2989 = _ctrlsignals_T_293 ? 2'h2 : _ctrlsignals_T_2988; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2990 = _ctrlsignals_T_291 ? 2'h1 : _ctrlsignals_T_2989; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2991 = _ctrlsignals_T_289 ? 2'h2 : _ctrlsignals_T_2990; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2992 = _ctrlsignals_T_287 ? 2'h1 : _ctrlsignals_T_2991; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2993 = _ctrlsignals_T_285 ? 2'h2 : _ctrlsignals_T_2992; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2994 = _ctrlsignals_T_283 ? 2'h1 : _ctrlsignals_T_2993; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2995 = _ctrlsignals_T_281 ? 2'h2 : _ctrlsignals_T_2994; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2996 = _ctrlsignals_T_279 ? 2'h3 : _ctrlsignals_T_2995; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2997 = _ctrlsignals_T_277 ? 2'h1 : _ctrlsignals_T_2996; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2998 = _ctrlsignals_T_275 ? 2'h2 : _ctrlsignals_T_2997; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_2999 = _ctrlsignals_T_273 ? 2'h3 : _ctrlsignals_T_2998; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3000 = _ctrlsignals_T_271 ? 2'h1 : _ctrlsignals_T_2999; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3001 = _ctrlsignals_T_269 ? 2'h2 : _ctrlsignals_T_3000; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3002 = _ctrlsignals_T_267 ? 2'h3 : _ctrlsignals_T_3001; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3003 = _ctrlsignals_T_265 ? 2'h1 : _ctrlsignals_T_3002; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3004 = _ctrlsignals_T_263 ? 2'h2 : _ctrlsignals_T_3003; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3005 = _ctrlsignals_T_261 ? 2'h3 : _ctrlsignals_T_3004; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3006 = _ctrlsignals_T_259 ? 2'h1 : _ctrlsignals_T_3005; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3007 = _ctrlsignals_T_257 ? 2'h2 : _ctrlsignals_T_3006; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3008 = _ctrlsignals_T_255 ? 2'h3 : _ctrlsignals_T_3007; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3009 = _ctrlsignals_T_253 ? 2'h1 : _ctrlsignals_T_3008; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3010 = _ctrlsignals_T_251 ? 2'h2 : _ctrlsignals_T_3009; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3011 = _ctrlsignals_T_249 ? 2'h1 : _ctrlsignals_T_3010; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3012 = _ctrlsignals_T_247 ? 2'h2 : _ctrlsignals_T_3011; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3013 = _ctrlsignals_T_245 ? 2'h1 : _ctrlsignals_T_3012; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3014 = _ctrlsignals_T_243 ? 2'h2 : _ctrlsignals_T_3013; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3015 = _ctrlsignals_T_241 ? 2'h3 : _ctrlsignals_T_3014; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3016 = _ctrlsignals_T_239 ? 2'h1 : _ctrlsignals_T_3015; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3017 = _ctrlsignals_T_237 ? 2'h1 : _ctrlsignals_T_3016; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3018 = _ctrlsignals_T_235 ? 2'h2 : _ctrlsignals_T_3017; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3019 = _ctrlsignals_T_233 ? 2'h1 : _ctrlsignals_T_3018; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3020 = _ctrlsignals_T_231 ? 2'h1 : _ctrlsignals_T_3019; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3021 = _ctrlsignals_T_229 ? 2'h2 : _ctrlsignals_T_3020; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3022 = _ctrlsignals_T_227 ? 2'h1 : _ctrlsignals_T_3021; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3023 = _ctrlsignals_T_225 ? 2'h2 : _ctrlsignals_T_3022; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3024 = _ctrlsignals_T_223 ? 2'h3 : _ctrlsignals_T_3023; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3025 = _ctrlsignals_T_221 ? 2'h1 : _ctrlsignals_T_3024; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3026 = _ctrlsignals_T_219 ? 2'h2 : _ctrlsignals_T_3025; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3027 = _ctrlsignals_T_217 ? 2'h1 : _ctrlsignals_T_3026; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3028 = _ctrlsignals_T_215 ? 2'h2 : _ctrlsignals_T_3027; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3029 = _ctrlsignals_T_213 ? 2'h1 : _ctrlsignals_T_3028; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3030 = _ctrlsignals_T_211 ? 2'h2 : _ctrlsignals_T_3029; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3031 = _ctrlsignals_T_209 ? 2'h1 : _ctrlsignals_T_3030; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3032 = _ctrlsignals_T_207 ? 2'h2 : _ctrlsignals_T_3031; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3033 = _ctrlsignals_T_205 ? 2'h1 : _ctrlsignals_T_3032; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3034 = _ctrlsignals_T_203 ? 2'h2 : _ctrlsignals_T_3033; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3035 = _ctrlsignals_T_201 ? 2'h1 : _ctrlsignals_T_3034; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3036 = _ctrlsignals_T_199 ? 2'h2 : _ctrlsignals_T_3035; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3037 = _ctrlsignals_T_197 ? 2'h1 : _ctrlsignals_T_3036; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3038 = _ctrlsignals_T_195 ? 2'h2 : _ctrlsignals_T_3037; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3039 = _ctrlsignals_T_193 ? 2'h1 : _ctrlsignals_T_3038; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3040 = _ctrlsignals_T_191 ? 2'h2 : _ctrlsignals_T_3039; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3041 = _ctrlsignals_T_189 ? 2'h1 : _ctrlsignals_T_3040; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3042 = _ctrlsignals_T_187 ? 2'h2 : _ctrlsignals_T_3041; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3043 = _ctrlsignals_T_185 ? 2'h1 : _ctrlsignals_T_3042; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3044 = _ctrlsignals_T_183 ? 2'h2 : _ctrlsignals_T_3043; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3045 = _ctrlsignals_T_181 ? 2'h1 : _ctrlsignals_T_3044; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3046 = _ctrlsignals_T_179 ? 2'h1 : _ctrlsignals_T_3045; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3047 = _ctrlsignals_T_177 ? 2'h1 : _ctrlsignals_T_3046; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3048 = _ctrlsignals_T_175 ? 2'h1 : _ctrlsignals_T_3047; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3049 = _ctrlsignals_T_173 ? 2'h1 : _ctrlsignals_T_3048; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3050 = _ctrlsignals_T_171 ? 2'h1 : _ctrlsignals_T_3049; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3051 = _ctrlsignals_T_169 ? 2'h1 : _ctrlsignals_T_3050; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3052 = _ctrlsignals_T_167 ? 2'h1 : _ctrlsignals_T_3051; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3053 = _ctrlsignals_T_165 ? 2'h1 : _ctrlsignals_T_3052; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3054 = _ctrlsignals_T_163 ? 2'h1 : _ctrlsignals_T_3053; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3055 = _ctrlsignals_T_161 ? 2'h1 : _ctrlsignals_T_3054; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3056 = _ctrlsignals_T_159 ? 2'h1 : _ctrlsignals_T_3055; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3057 = _ctrlsignals_T_143 ? 2'h1 : _ctrlsignals_T_3056; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3058 = _ctrlsignals_T_155 ? 2'h1 : _ctrlsignals_T_3057; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3059 = _ctrlsignals_T_153 ? 2'h1 : _ctrlsignals_T_3058; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3060 = _ctrlsignals_T_151 ? 2'h1 : _ctrlsignals_T_3059; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3061 = _ctrlsignals_T_149 ? 2'h1 : _ctrlsignals_T_3060; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3062 = _ctrlsignals_T_147 ? 2'h1 : _ctrlsignals_T_3061; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3063 = _ctrlsignals_T_145 ? 2'h1 : _ctrlsignals_T_3062; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3064 = _ctrlsignals_T_143 ? 2'h1 : _ctrlsignals_T_3063; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3065 = _ctrlsignals_T_141 ? 2'h1 : _ctrlsignals_T_3064; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3066 = _ctrlsignals_T_139 ? 2'h1 : _ctrlsignals_T_3065; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3067 = _ctrlsignals_T_137 ? 2'h1 : _ctrlsignals_T_3066; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3068 = _ctrlsignals_T_135 ? 2'h1 : _ctrlsignals_T_3067; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3069 = _ctrlsignals_T_133 ? 2'h1 : _ctrlsignals_T_3068; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3070 = _ctrlsignals_T_131 ? 2'h1 : _ctrlsignals_T_3069; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3071 = _ctrlsignals_T_129 ? 2'h1 : _ctrlsignals_T_3070; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3072 = _ctrlsignals_T_127 ? 2'h1 : _ctrlsignals_T_3071; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3073 = _ctrlsignals_T_125 ? 2'h1 : _ctrlsignals_T_3072; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3074 = _ctrlsignals_T_123 ? 2'h1 : _ctrlsignals_T_3073; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3075 = _ctrlsignals_T_121 ? 2'h1 : _ctrlsignals_T_3074; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3076 = _ctrlsignals_T_119 ? 2'h1 : _ctrlsignals_T_3075; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3077 = _ctrlsignals_T_117 ? 2'h1 : _ctrlsignals_T_3076; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3078 = _ctrlsignals_T_115 ? 2'h1 : _ctrlsignals_T_3077; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3079 = _ctrlsignals_T_113 ? 2'h1 : _ctrlsignals_T_3078; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3080 = _ctrlsignals_T_111 ? 2'h1 : _ctrlsignals_T_3079; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3081 = _ctrlsignals_T_109 ? 2'h1 : _ctrlsignals_T_3080; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3082 = _ctrlsignals_T_107 ? 2'h1 : _ctrlsignals_T_3081; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3083 = _ctrlsignals_T_105 ? 2'h1 : _ctrlsignals_T_3082; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3084 = _ctrlsignals_T_103 ? 2'h1 : _ctrlsignals_T_3083; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3085 = _ctrlsignals_T_101 ? 2'h1 : _ctrlsignals_T_3084; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3086 = _ctrlsignals_T_99 ? 2'h1 : _ctrlsignals_T_3085; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3087 = _ctrlsignals_T_97 ? 2'h1 : _ctrlsignals_T_3086; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3088 = _ctrlsignals_T_95 ? 2'h1 : _ctrlsignals_T_3087; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3089 = _ctrlsignals_T_93 ? 2'h1 : _ctrlsignals_T_3088; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3090 = _ctrlsignals_T_91 ? 2'h1 : _ctrlsignals_T_3089; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3091 = _ctrlsignals_T_89 ? 2'h1 : _ctrlsignals_T_3090; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3092 = _ctrlsignals_T_87 ? 2'h1 : _ctrlsignals_T_3091; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3093 = _ctrlsignals_T_85 ? 2'h1 : _ctrlsignals_T_3092; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3094 = _ctrlsignals_T_83 ? 2'h1 : _ctrlsignals_T_3093; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3095 = _ctrlsignals_T_81 ? 2'h1 : _ctrlsignals_T_3094; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3096 = _ctrlsignals_T_79 ? 2'h1 : _ctrlsignals_T_3095; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3097 = _ctrlsignals_T_77 ? 2'h1 : _ctrlsignals_T_3096; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3098 = _ctrlsignals_T_75 ? 2'h1 : _ctrlsignals_T_3097; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3099 = _ctrlsignals_T_73 ? 2'h1 : _ctrlsignals_T_3098; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3100 = _ctrlsignals_T_71 ? 2'h1 : _ctrlsignals_T_3099; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3101 = _ctrlsignals_T_69 ? 2'h1 : _ctrlsignals_T_3100; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3102 = _ctrlsignals_T_67 ? 2'h1 : _ctrlsignals_T_3101; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3103 = _ctrlsignals_T_65 ? 2'h1 : _ctrlsignals_T_3102; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3104 = _ctrlsignals_T_63 ? 2'h1 : _ctrlsignals_T_3103; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3105 = _ctrlsignals_T_61 ? 2'h1 : _ctrlsignals_T_3104; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3106 = _ctrlsignals_T_59 ? 2'h1 : _ctrlsignals_T_3105; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3107 = _ctrlsignals_T_57 ? 2'h1 : _ctrlsignals_T_3106; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3108 = _ctrlsignals_T_55 ? 2'h1 : _ctrlsignals_T_3107; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3109 = _ctrlsignals_T_53 ? 2'h1 : _ctrlsignals_T_3108; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3110 = _ctrlsignals_T_51 ? 2'h1 : _ctrlsignals_T_3109; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3111 = _ctrlsignals_T_49 ? 2'h1 : _ctrlsignals_T_3110; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3112 = _ctrlsignals_T_47 ? 2'h3 : _ctrlsignals_T_3111; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3113 = _ctrlsignals_T_45 ? 2'h3 : _ctrlsignals_T_3112; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3114 = _ctrlsignals_T_43 ? 2'h3 : _ctrlsignals_T_3113; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3115 = _ctrlsignals_T_41 ? 2'h1 : _ctrlsignals_T_3114; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3116 = _ctrlsignals_T_39 ? 2'h1 : _ctrlsignals_T_3115; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3117 = _ctrlsignals_T_37 ? 2'h1 : _ctrlsignals_T_3116; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3118 = _ctrlsignals_T_35 ? 2'h0 : _ctrlsignals_T_3117; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3119 = _ctrlsignals_T_33 ? 2'h0 : _ctrlsignals_T_3118; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3120 = _ctrlsignals_T_31 ? 2'h0 : _ctrlsignals_T_3119; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3121 = _ctrlsignals_T_29 ? 2'h1 : _ctrlsignals_T_3120; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3122 = _ctrlsignals_T_27 ? 2'h1 : _ctrlsignals_T_3121; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3123 = _ctrlsignals_T_25 ? 2'h1 : _ctrlsignals_T_3122; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3124 = _ctrlsignals_T_23 ? 2'h1 : _ctrlsignals_T_3123; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3125 = _ctrlsignals_T_21 ? 2'h1 : _ctrlsignals_T_3124; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3126 = _ctrlsignals_T_19 ? 2'h1 : _ctrlsignals_T_3125; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3127 = _ctrlsignals_T_17 ? 2'h1 : _ctrlsignals_T_3126; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3128 = _ctrlsignals_T_15 ? 2'h3 : _ctrlsignals_T_3127; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3129 = _ctrlsignals_T_13 ? 2'h1 : _ctrlsignals_T_3128; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3130 = _ctrlsignals_T_11 ? 2'h2 : _ctrlsignals_T_3129; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3131 = _ctrlsignals_T_9 ? 2'h2 : _ctrlsignals_T_3130; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3132 = _ctrlsignals_T_7 ? 2'h2 : _ctrlsignals_T_3131; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3133 = _ctrlsignals_T_5 ? 2'h2 : _ctrlsignals_T_3132; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_3134 = _ctrlsignals_T_3 ? 2'h2 : _ctrlsignals_T_3133; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3136 = _ctrlsignals_T_481 ? 3'h7 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3137 = _ctrlsignals_T_479 ? 3'h0 : _ctrlsignals_T_3136; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3138 = _ctrlsignals_T_477 ? 3'h0 : _ctrlsignals_T_3137; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3139 = _ctrlsignals_T_475 ? 3'h0 : _ctrlsignals_T_3138; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3140 = _ctrlsignals_T_473 ? 3'h6 : _ctrlsignals_T_3139; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3141 = _ctrlsignals_T_471 ? 3'h0 : _ctrlsignals_T_3140; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3142 = _ctrlsignals_T_469 ? 3'h0 : _ctrlsignals_T_3141; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3143 = _ctrlsignals_T_467 ? 3'h0 : _ctrlsignals_T_3142; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3144 = _ctrlsignals_T_465 ? 3'h0 : _ctrlsignals_T_3143; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3145 = _ctrlsignals_T_463 ? 3'h0 : _ctrlsignals_T_3144; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3146 = _ctrlsignals_T_461 ? 3'h0 : _ctrlsignals_T_3145; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3147 = _ctrlsignals_T_459 ? 3'h0 : _ctrlsignals_T_3146; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3148 = _ctrlsignals_T_445 ? 3'h0 : _ctrlsignals_T_3147; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3149 = _ctrlsignals_T_443 ? 3'h0 : _ctrlsignals_T_3148; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3150 = _ctrlsignals_T_453 ? 3'h0 : _ctrlsignals_T_3149; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3151 = _ctrlsignals_T_451 ? 3'h0 : _ctrlsignals_T_3150; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3152 = _ctrlsignals_T_449 ? 3'h0 : _ctrlsignals_T_3151; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3153 = _ctrlsignals_T_447 ? 3'h0 : _ctrlsignals_T_3152; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3154 = _ctrlsignals_T_445 ? 3'h0 : _ctrlsignals_T_3153; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3155 = _ctrlsignals_T_443 ? 3'h0 : _ctrlsignals_T_3154; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3156 = _ctrlsignals_T_441 ? 3'h0 : _ctrlsignals_T_3155; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3157 = _ctrlsignals_T_439 ? 3'h0 : _ctrlsignals_T_3156; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3158 = _ctrlsignals_T_437 ? 3'h0 : _ctrlsignals_T_3157; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3159 = _ctrlsignals_T_435 ? 3'h0 : _ctrlsignals_T_3158; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3160 = _ctrlsignals_T_433 ? 3'h0 : _ctrlsignals_T_3159; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3161 = _ctrlsignals_T_431 ? 3'h0 : _ctrlsignals_T_3160; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3162 = _ctrlsignals_T_429 ? 3'h0 : _ctrlsignals_T_3161; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3163 = _ctrlsignals_T_427 ? 3'h0 : _ctrlsignals_T_3162; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3164 = _ctrlsignals_T_425 ? 3'h0 : _ctrlsignals_T_3163; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3165 = _ctrlsignals_T_423 ? 3'h0 : _ctrlsignals_T_3164; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3166 = _ctrlsignals_T_421 ? 3'h0 : _ctrlsignals_T_3165; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3167 = _ctrlsignals_T_419 ? 3'h0 : _ctrlsignals_T_3166; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3168 = _ctrlsignals_T_417 ? 3'h0 : _ctrlsignals_T_3167; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3169 = _ctrlsignals_T_415 ? 3'h0 : _ctrlsignals_T_3168; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3170 = _ctrlsignals_T_413 ? 3'h0 : _ctrlsignals_T_3169; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3171 = _ctrlsignals_T_411 ? 3'h0 : _ctrlsignals_T_3170; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3172 = _ctrlsignals_T_409 ? 3'h0 : _ctrlsignals_T_3171; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3173 = _ctrlsignals_T_407 ? 3'h0 : _ctrlsignals_T_3172; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3174 = _ctrlsignals_T_405 ? 3'h0 : _ctrlsignals_T_3173; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3175 = _ctrlsignals_T_403 ? 3'h0 : _ctrlsignals_T_3174; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3176 = _ctrlsignals_T_401 ? 3'h0 : _ctrlsignals_T_3175; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3177 = _ctrlsignals_T_399 ? 3'h0 : _ctrlsignals_T_3176; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3178 = _ctrlsignals_T_397 ? 3'h0 : _ctrlsignals_T_3177; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3179 = _ctrlsignals_T_395 ? 3'h0 : _ctrlsignals_T_3178; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3180 = _ctrlsignals_T_393 ? 3'h0 : _ctrlsignals_T_3179; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3181 = _ctrlsignals_T_391 ? 3'h0 : _ctrlsignals_T_3180; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3182 = _ctrlsignals_T_389 ? 3'h0 : _ctrlsignals_T_3181; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3183 = _ctrlsignals_T_387 ? 3'h0 : _ctrlsignals_T_3182; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3184 = _ctrlsignals_T_385 ? 3'h0 : _ctrlsignals_T_3183; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3185 = _ctrlsignals_T_383 ? 3'h0 : _ctrlsignals_T_3184; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3186 = _ctrlsignals_T_381 ? 3'h0 : _ctrlsignals_T_3185; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3187 = _ctrlsignals_T_379 ? 3'h0 : _ctrlsignals_T_3186; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3188 = _ctrlsignals_T_377 ? 3'h0 : _ctrlsignals_T_3187; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3189 = _ctrlsignals_T_375 ? 3'h0 : _ctrlsignals_T_3188; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3190 = _ctrlsignals_T_373 ? 3'h0 : _ctrlsignals_T_3189; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3191 = _ctrlsignals_T_371 ? 3'h0 : _ctrlsignals_T_3190; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3192 = _ctrlsignals_T_369 ? 3'h6 : _ctrlsignals_T_3191; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3193 = _ctrlsignals_T_367 ? 3'h0 : _ctrlsignals_T_3192; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3194 = _ctrlsignals_T_365 ? 3'h0 : _ctrlsignals_T_3193; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3195 = _ctrlsignals_T_363 ? 3'h0 : _ctrlsignals_T_3194; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3196 = _ctrlsignals_T_361 ? 3'h0 : _ctrlsignals_T_3195; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3197 = _ctrlsignals_T_359 ? 3'h0 : _ctrlsignals_T_3196; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3198 = _ctrlsignals_T_357 ? 3'h0 : _ctrlsignals_T_3197; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3199 = _ctrlsignals_T_355 ? 3'h0 : _ctrlsignals_T_3198; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3200 = _ctrlsignals_T_353 ? 3'h0 : _ctrlsignals_T_3199; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3201 = _ctrlsignals_T_351 ? 3'h0 : _ctrlsignals_T_3200; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3202 = _ctrlsignals_T_349 ? 3'h0 : _ctrlsignals_T_3201; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3203 = _ctrlsignals_T_347 ? 3'h0 : _ctrlsignals_T_3202; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3204 = _ctrlsignals_T_345 ? 3'h0 : _ctrlsignals_T_3203; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3205 = _ctrlsignals_T_343 ? 3'h6 : _ctrlsignals_T_3204; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3206 = _ctrlsignals_T_341 ? 3'h0 : _ctrlsignals_T_3205; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3207 = _ctrlsignals_T_339 ? 3'h7 : _ctrlsignals_T_3206; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3208 = _ctrlsignals_T_337 ? 3'h0 : _ctrlsignals_T_3207; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3209 = _ctrlsignals_T_335 ? 3'h6 : _ctrlsignals_T_3208; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3210 = _ctrlsignals_T_333 ? 3'h0 : _ctrlsignals_T_3209; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3211 = _ctrlsignals_T_331 ? 3'h0 : _ctrlsignals_T_3210; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3212 = _ctrlsignals_T_329 ? 3'h7 : _ctrlsignals_T_3211; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3213 = _ctrlsignals_T_327 ? 3'h0 : _ctrlsignals_T_3212; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3214 = _ctrlsignals_T_325 ? 3'h6 : _ctrlsignals_T_3213; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3215 = _ctrlsignals_T_323 ? 3'h0 : _ctrlsignals_T_3214; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3216 = _ctrlsignals_T_321 ? 3'h0 : _ctrlsignals_T_3215; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3217 = _ctrlsignals_T_319 ? 3'h6 : _ctrlsignals_T_3216; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3218 = _ctrlsignals_T_317 ? 3'h0 : _ctrlsignals_T_3217; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3219 = _ctrlsignals_T_315 ? 3'h0 : _ctrlsignals_T_3218; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3220 = _ctrlsignals_T_313 ? 3'h6 : _ctrlsignals_T_3219; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3221 = _ctrlsignals_T_311 ? 3'h0 : _ctrlsignals_T_3220; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3222 = _ctrlsignals_T_309 ? 3'h0 : _ctrlsignals_T_3221; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3223 = _ctrlsignals_T_307 ? 3'h0 : _ctrlsignals_T_3222; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3224 = _ctrlsignals_T_305 ? 3'h0 : _ctrlsignals_T_3223; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3225 = _ctrlsignals_T_303 ? 3'h0 : _ctrlsignals_T_3224; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3226 = _ctrlsignals_T_301 ? 3'h0 : _ctrlsignals_T_3225; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3227 = _ctrlsignals_T_299 ? 3'h0 : _ctrlsignals_T_3226; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3228 = _ctrlsignals_T_297 ? 3'h0 : _ctrlsignals_T_3227; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3229 = _ctrlsignals_T_295 ? 3'h0 : _ctrlsignals_T_3228; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3230 = _ctrlsignals_T_293 ? 3'h0 : _ctrlsignals_T_3229; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3231 = _ctrlsignals_T_291 ? 3'h0 : _ctrlsignals_T_3230; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3232 = _ctrlsignals_T_289 ? 3'h0 : _ctrlsignals_T_3231; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3233 = _ctrlsignals_T_287 ? 3'h0 : _ctrlsignals_T_3232; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3234 = _ctrlsignals_T_285 ? 3'h0 : _ctrlsignals_T_3233; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3235 = _ctrlsignals_T_283 ? 3'h0 : _ctrlsignals_T_3234; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3236 = _ctrlsignals_T_281 ? 3'h0 : _ctrlsignals_T_3235; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3237 = _ctrlsignals_T_279 ? 3'h6 : _ctrlsignals_T_3236; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3238 = _ctrlsignals_T_277 ? 3'h0 : _ctrlsignals_T_3237; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3239 = _ctrlsignals_T_275 ? 3'h0 : _ctrlsignals_T_3238; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3240 = _ctrlsignals_T_273 ? 3'h6 : _ctrlsignals_T_3239; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3241 = _ctrlsignals_T_271 ? 3'h0 : _ctrlsignals_T_3240; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3242 = _ctrlsignals_T_269 ? 3'h0 : _ctrlsignals_T_3241; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3243 = _ctrlsignals_T_267 ? 3'h6 : _ctrlsignals_T_3242; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3244 = _ctrlsignals_T_265 ? 3'h0 : _ctrlsignals_T_3243; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3245 = _ctrlsignals_T_263 ? 3'h0 : _ctrlsignals_T_3244; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3246 = _ctrlsignals_T_261 ? 3'h6 : _ctrlsignals_T_3245; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3247 = _ctrlsignals_T_259 ? 3'h0 : _ctrlsignals_T_3246; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3248 = _ctrlsignals_T_257 ? 3'h0 : _ctrlsignals_T_3247; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3249 = _ctrlsignals_T_255 ? 3'h6 : _ctrlsignals_T_3248; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3250 = _ctrlsignals_T_253 ? 3'h0 : _ctrlsignals_T_3249; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3251 = _ctrlsignals_T_251 ? 3'h0 : _ctrlsignals_T_3250; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3252 = _ctrlsignals_T_249 ? 3'h0 : _ctrlsignals_T_3251; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3253 = _ctrlsignals_T_247 ? 3'h0 : _ctrlsignals_T_3252; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3254 = _ctrlsignals_T_245 ? 3'h0 : _ctrlsignals_T_3253; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3255 = _ctrlsignals_T_243 ? 3'h0 : _ctrlsignals_T_3254; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3256 = _ctrlsignals_T_241 ? 3'h6 : _ctrlsignals_T_3255; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3257 = _ctrlsignals_T_239 ? 3'h0 : _ctrlsignals_T_3256; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3258 = _ctrlsignals_T_237 ? 3'h0 : _ctrlsignals_T_3257; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3259 = _ctrlsignals_T_235 ? 3'h0 : _ctrlsignals_T_3258; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3260 = _ctrlsignals_T_233 ? 3'h0 : _ctrlsignals_T_3259; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3261 = _ctrlsignals_T_231 ? 3'h0 : _ctrlsignals_T_3260; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3262 = _ctrlsignals_T_229 ? 3'h0 : _ctrlsignals_T_3261; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3263 = _ctrlsignals_T_227 ? 3'h0 : _ctrlsignals_T_3262; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3264 = _ctrlsignals_T_225 ? 3'h0 : _ctrlsignals_T_3263; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3265 = _ctrlsignals_T_223 ? 3'h6 : _ctrlsignals_T_3264; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3266 = _ctrlsignals_T_221 ? 3'h0 : _ctrlsignals_T_3265; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3267 = _ctrlsignals_T_219 ? 3'h0 : _ctrlsignals_T_3266; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3268 = _ctrlsignals_T_217 ? 3'h0 : _ctrlsignals_T_3267; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3269 = _ctrlsignals_T_215 ? 3'h0 : _ctrlsignals_T_3268; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3270 = _ctrlsignals_T_213 ? 3'h0 : _ctrlsignals_T_3269; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3271 = _ctrlsignals_T_211 ? 3'h0 : _ctrlsignals_T_3270; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3272 = _ctrlsignals_T_209 ? 3'h0 : _ctrlsignals_T_3271; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3273 = _ctrlsignals_T_207 ? 3'h0 : _ctrlsignals_T_3272; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3274 = _ctrlsignals_T_205 ? 3'h0 : _ctrlsignals_T_3273; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3275 = _ctrlsignals_T_203 ? 3'h0 : _ctrlsignals_T_3274; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3276 = _ctrlsignals_T_201 ? 3'h0 : _ctrlsignals_T_3275; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3277 = _ctrlsignals_T_199 ? 3'h0 : _ctrlsignals_T_3276; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3278 = _ctrlsignals_T_197 ? 3'h0 : _ctrlsignals_T_3277; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3279 = _ctrlsignals_T_195 ? 3'h0 : _ctrlsignals_T_3278; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3280 = _ctrlsignals_T_193 ? 3'h0 : _ctrlsignals_T_3279; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3281 = _ctrlsignals_T_191 ? 3'h0 : _ctrlsignals_T_3280; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3282 = _ctrlsignals_T_189 ? 3'h0 : _ctrlsignals_T_3281; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3283 = _ctrlsignals_T_187 ? 3'h0 : _ctrlsignals_T_3282; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3284 = _ctrlsignals_T_185 ? 3'h0 : _ctrlsignals_T_3283; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3285 = _ctrlsignals_T_183 ? 3'h0 : _ctrlsignals_T_3284; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3286 = _ctrlsignals_T_181 ? 3'h0 : _ctrlsignals_T_3285; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3287 = _ctrlsignals_T_179 ? 3'h0 : _ctrlsignals_T_3286; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3288 = _ctrlsignals_T_177 ? 3'h0 : _ctrlsignals_T_3287; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3289 = _ctrlsignals_T_175 ? 3'h0 : _ctrlsignals_T_3288; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3290 = _ctrlsignals_T_173 ? 3'h0 : _ctrlsignals_T_3289; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3291 = _ctrlsignals_T_171 ? 3'h0 : _ctrlsignals_T_3290; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3292 = _ctrlsignals_T_169 ? 3'h0 : _ctrlsignals_T_3291; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3293 = _ctrlsignals_T_167 ? 3'h0 : _ctrlsignals_T_3292; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3294 = _ctrlsignals_T_165 ? 3'h0 : _ctrlsignals_T_3293; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3295 = _ctrlsignals_T_163 ? 3'h0 : _ctrlsignals_T_3294; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3296 = _ctrlsignals_T_161 ? 3'h0 : _ctrlsignals_T_3295; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3297 = _ctrlsignals_T_159 ? 3'h0 : _ctrlsignals_T_3296; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3298 = _ctrlsignals_T_143 ? 3'h0 : _ctrlsignals_T_3297; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3299 = _ctrlsignals_T_155 ? 3'h0 : _ctrlsignals_T_3298; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3300 = _ctrlsignals_T_153 ? 3'h0 : _ctrlsignals_T_3299; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3301 = _ctrlsignals_T_151 ? 3'h0 : _ctrlsignals_T_3300; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3302 = _ctrlsignals_T_149 ? 3'h0 : _ctrlsignals_T_3301; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3303 = _ctrlsignals_T_147 ? 3'h0 : _ctrlsignals_T_3302; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3304 = _ctrlsignals_T_145 ? 3'h0 : _ctrlsignals_T_3303; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3305 = _ctrlsignals_T_143 ? 3'h0 : _ctrlsignals_T_3304; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3306 = _ctrlsignals_T_141 ? 3'h0 : _ctrlsignals_T_3305; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3307 = _ctrlsignals_T_139 ? 3'h0 : _ctrlsignals_T_3306; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3308 = _ctrlsignals_T_137 ? 3'h0 : _ctrlsignals_T_3307; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3309 = _ctrlsignals_T_135 ? 3'h0 : _ctrlsignals_T_3308; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3310 = _ctrlsignals_T_133 ? 3'h0 : _ctrlsignals_T_3309; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3311 = _ctrlsignals_T_131 ? 3'h0 : _ctrlsignals_T_3310; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3312 = _ctrlsignals_T_129 ? 3'h0 : _ctrlsignals_T_3311; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3313 = _ctrlsignals_T_127 ? 3'h0 : _ctrlsignals_T_3312; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3314 = _ctrlsignals_T_125 ? 3'h0 : _ctrlsignals_T_3313; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3315 = _ctrlsignals_T_123 ? 3'h0 : _ctrlsignals_T_3314; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3316 = _ctrlsignals_T_121 ? 3'h0 : _ctrlsignals_T_3315; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3317 = _ctrlsignals_T_119 ? 3'h0 : _ctrlsignals_T_3316; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3318 = _ctrlsignals_T_117 ? 3'h0 : _ctrlsignals_T_3317; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3319 = _ctrlsignals_T_115 ? 3'h0 : _ctrlsignals_T_3318; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3320 = _ctrlsignals_T_113 ? 3'h0 : _ctrlsignals_T_3319; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3321 = _ctrlsignals_T_111 ? 3'h0 : _ctrlsignals_T_3320; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3322 = _ctrlsignals_T_109 ? 3'h0 : _ctrlsignals_T_3321; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3323 = _ctrlsignals_T_107 ? 3'h0 : _ctrlsignals_T_3322; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3324 = _ctrlsignals_T_105 ? 3'h4 : _ctrlsignals_T_3323; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3325 = _ctrlsignals_T_103 ? 3'h4 : _ctrlsignals_T_3324; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3326 = _ctrlsignals_T_101 ? 3'h4 : _ctrlsignals_T_3325; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3327 = _ctrlsignals_T_99 ? 3'h0 : _ctrlsignals_T_3326; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3328 = _ctrlsignals_T_97 ? 3'h0 : _ctrlsignals_T_3327; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3329 = _ctrlsignals_T_95 ? 3'h0 : _ctrlsignals_T_3328; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3330 = _ctrlsignals_T_93 ? 3'h0 : _ctrlsignals_T_3329; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3331 = _ctrlsignals_T_91 ? 3'h0 : _ctrlsignals_T_3330; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3332 = _ctrlsignals_T_89 ? 3'h0 : _ctrlsignals_T_3331; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3333 = _ctrlsignals_T_87 ? 3'h0 : _ctrlsignals_T_3332; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3334 = _ctrlsignals_T_85 ? 3'h0 : _ctrlsignals_T_3333; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3335 = _ctrlsignals_T_83 ? 3'h0 : _ctrlsignals_T_3334; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3336 = _ctrlsignals_T_81 ? 3'h0 : _ctrlsignals_T_3335; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3337 = _ctrlsignals_T_79 ? 3'h0 : _ctrlsignals_T_3336; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3338 = _ctrlsignals_T_77 ? 3'h0 : _ctrlsignals_T_3337; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3339 = _ctrlsignals_T_75 ? 3'h0 : _ctrlsignals_T_3338; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3340 = _ctrlsignals_T_73 ? 3'h0 : _ctrlsignals_T_3339; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3341 = _ctrlsignals_T_71 ? 3'h0 : _ctrlsignals_T_3340; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3342 = _ctrlsignals_T_69 ? 3'h0 : _ctrlsignals_T_3341; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3343 = _ctrlsignals_T_67 ? 3'h3 : _ctrlsignals_T_3342; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3344 = _ctrlsignals_T_65 ? 3'h1 : _ctrlsignals_T_3343; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3345 = _ctrlsignals_T_63 ? 3'h1 : _ctrlsignals_T_3344; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3346 = _ctrlsignals_T_61 ? 3'h1 : _ctrlsignals_T_3345; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3347 = _ctrlsignals_T_59 ? 3'h0 : _ctrlsignals_T_3346; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3348 = _ctrlsignals_T_57 ? 3'h0 : _ctrlsignals_T_3347; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3349 = _ctrlsignals_T_55 ? 3'h0 : _ctrlsignals_T_3348; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3350 = _ctrlsignals_T_53 ? 3'h0 : _ctrlsignals_T_3349; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3351 = _ctrlsignals_T_51 ? 3'h0 : _ctrlsignals_T_3350; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3352 = _ctrlsignals_T_49 ? 3'h0 : _ctrlsignals_T_3351; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3353 = _ctrlsignals_T_47 ? 3'h7 : _ctrlsignals_T_3352; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3354 = _ctrlsignals_T_45 ? 3'h7 : _ctrlsignals_T_3353; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3355 = _ctrlsignals_T_43 ? 3'h7 : _ctrlsignals_T_3354; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3356 = _ctrlsignals_T_41 ? 3'h0 : _ctrlsignals_T_3355; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3357 = _ctrlsignals_T_39 ? 3'h0 : _ctrlsignals_T_3356; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3358 = _ctrlsignals_T_37 ? 3'h0 : _ctrlsignals_T_3357; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3359 = _ctrlsignals_T_35 ? 3'h3 : _ctrlsignals_T_3358; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3360 = _ctrlsignals_T_33 ? 3'h0 : _ctrlsignals_T_3359; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3361 = _ctrlsignals_T_31 ? 3'h5 : _ctrlsignals_T_3360; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3362 = _ctrlsignals_T_29 ? 3'h2 : _ctrlsignals_T_3361; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3363 = _ctrlsignals_T_27 ? 3'h2 : _ctrlsignals_T_3362; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3364 = _ctrlsignals_T_25 ? 3'h2 : _ctrlsignals_T_3363; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3365 = _ctrlsignals_T_23 ? 3'h2 : _ctrlsignals_T_3364; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3366 = _ctrlsignals_T_21 ? 3'h2 : _ctrlsignals_T_3365; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3367 = _ctrlsignals_T_19 ? 3'h2 : _ctrlsignals_T_3366; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3368 = _ctrlsignals_T_17 ? 3'h0 : _ctrlsignals_T_3367; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3369 = _ctrlsignals_T_15 ? 3'h7 : _ctrlsignals_T_3368; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3370 = _ctrlsignals_T_13 ? 3'h2 : _ctrlsignals_T_3369; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3371 = _ctrlsignals_T_11 ? 3'h2 : _ctrlsignals_T_3370; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3372 = _ctrlsignals_T_9 ? 3'h2 : _ctrlsignals_T_3371; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3373 = _ctrlsignals_T_7 ? 3'h2 : _ctrlsignals_T_3372; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3374 = _ctrlsignals_T_5 ? 3'h2 : _ctrlsignals_T_3373; // @[Lookup.scala 34:39]
  wire [2:0] _ctrlsignals_T_3375 = _ctrlsignals_T_3 ? 3'h2 : _ctrlsignals_T_3374; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3617 = _ctrlsignals_T_483 ? 6'h0 : 6'h3f; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3618 = _ctrlsignals_T_481 ? 6'h0 : _ctrlsignals_T_3617; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3619 = _ctrlsignals_T_479 ? 6'h0 : _ctrlsignals_T_3618; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3620 = _ctrlsignals_T_477 ? 6'h0 : _ctrlsignals_T_3619; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3621 = _ctrlsignals_T_475 ? 6'h0 : _ctrlsignals_T_3620; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3622 = _ctrlsignals_T_473 ? 6'h0 : _ctrlsignals_T_3621; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3623 = _ctrlsignals_T_471 ? 6'h0 : _ctrlsignals_T_3622; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3624 = _ctrlsignals_T_469 ? 6'h0 : _ctrlsignals_T_3623; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3625 = _ctrlsignals_T_467 ? 6'h12 : _ctrlsignals_T_3624; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3626 = _ctrlsignals_T_465 ? 6'h20 : _ctrlsignals_T_3625; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3627 = _ctrlsignals_T_463 ? 6'h21 : _ctrlsignals_T_3626; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3628 = _ctrlsignals_T_461 ? 6'h18 : _ctrlsignals_T_3627; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3629 = _ctrlsignals_T_459 ? 6'h19 : _ctrlsignals_T_3628; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3630 = _ctrlsignals_T_445 ? 6'h16 : _ctrlsignals_T_3629; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3631 = _ctrlsignals_T_443 ? 6'h16 : _ctrlsignals_T_3630; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3632 = _ctrlsignals_T_453 ? 6'h14 : _ctrlsignals_T_3631; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3633 = _ctrlsignals_T_451 ? 6'h14 : _ctrlsignals_T_3632; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3634 = _ctrlsignals_T_449 ? 6'h15 : _ctrlsignals_T_3633; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3635 = _ctrlsignals_T_447 ? 6'h15 : _ctrlsignals_T_3634; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3636 = _ctrlsignals_T_445 ? 6'h16 : _ctrlsignals_T_3635; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3637 = _ctrlsignals_T_443 ? 6'h16 : _ctrlsignals_T_3636; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3638 = _ctrlsignals_T_441 ? 6'h10 : _ctrlsignals_T_3637; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3639 = _ctrlsignals_T_439 ? 6'h11 : _ctrlsignals_T_3638; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3640 = _ctrlsignals_T_437 ? 6'h12 : _ctrlsignals_T_3639; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3641 = _ctrlsignals_T_435 ? 6'h13 : _ctrlsignals_T_3640; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3642 = _ctrlsignals_T_433 ? 6'h10 : _ctrlsignals_T_3641; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3643 = _ctrlsignals_T_431 ? 6'h11 : _ctrlsignals_T_3642; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3644 = _ctrlsignals_T_429 ? 6'h12 : _ctrlsignals_T_3643; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3645 = _ctrlsignals_T_427 ? 6'h13 : _ctrlsignals_T_3644; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3646 = _ctrlsignals_T_425 ? 6'h1 : _ctrlsignals_T_3645; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3647 = _ctrlsignals_T_423 ? 6'h0 : _ctrlsignals_T_3646; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3648 = _ctrlsignals_T_421 ? 6'h0 : _ctrlsignals_T_3647; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3649 = _ctrlsignals_T_419 ? 6'h0 : _ctrlsignals_T_3648; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3650 = _ctrlsignals_T_417 ? 6'h2 : _ctrlsignals_T_3649; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3651 = _ctrlsignals_T_415 ? 6'h2 : _ctrlsignals_T_3650; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3652 = _ctrlsignals_T_413 ? 6'h0 : _ctrlsignals_T_3651; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3653 = _ctrlsignals_T_411 ? 6'h0 : _ctrlsignals_T_3652; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3654 = _ctrlsignals_T_409 ? 6'h3 : _ctrlsignals_T_3653; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3655 = _ctrlsignals_T_407 ? 6'h3 : _ctrlsignals_T_3654; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3656 = _ctrlsignals_T_405 ? 6'h1 : _ctrlsignals_T_3655; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3657 = _ctrlsignals_T_403 ? 6'h1 : _ctrlsignals_T_3656; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3658 = _ctrlsignals_T_401 ? 6'h1b : _ctrlsignals_T_3657; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3659 = _ctrlsignals_T_399 ? 6'h1b : _ctrlsignals_T_3658; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3660 = _ctrlsignals_T_397 ? 6'h1a : _ctrlsignals_T_3659; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3661 = _ctrlsignals_T_395 ? 6'h1a : _ctrlsignals_T_3660; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3662 = _ctrlsignals_T_393 ? 6'h19 : _ctrlsignals_T_3661; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3663 = _ctrlsignals_T_391 ? 6'h19 : _ctrlsignals_T_3662; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3664 = _ctrlsignals_T_389 ? 6'h18 : _ctrlsignals_T_3663; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3665 = _ctrlsignals_T_387 ? 6'h18 : _ctrlsignals_T_3664; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3666 = _ctrlsignals_T_385 ? 6'h17 : _ctrlsignals_T_3665; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3667 = _ctrlsignals_T_383 ? 6'h17 : _ctrlsignals_T_3666; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3668 = _ctrlsignals_T_381 ? 6'h16 : _ctrlsignals_T_3667; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3669 = _ctrlsignals_T_379 ? 6'h16 : _ctrlsignals_T_3668; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3670 = _ctrlsignals_T_377 ? 6'h15 : _ctrlsignals_T_3669; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3671 = _ctrlsignals_T_375 ? 6'h15 : _ctrlsignals_T_3670; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3672 = _ctrlsignals_T_373 ? 6'h14 : _ctrlsignals_T_3671; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3673 = _ctrlsignals_T_371 ? 6'h14 : _ctrlsignals_T_3672; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3674 = _ctrlsignals_T_369 ? 6'h13 : _ctrlsignals_T_3673; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3675 = _ctrlsignals_T_367 ? 6'h13 : _ctrlsignals_T_3674; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3676 = _ctrlsignals_T_365 ? 6'h13 : _ctrlsignals_T_3675; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3677 = _ctrlsignals_T_363 ? 6'h19 : _ctrlsignals_T_3676; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3678 = _ctrlsignals_T_361 ? 6'h18 : _ctrlsignals_T_3677; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3679 = _ctrlsignals_T_359 ? 6'h16 : _ctrlsignals_T_3678; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3680 = _ctrlsignals_T_357 ? 6'h17 : _ctrlsignals_T_3679; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3681 = _ctrlsignals_T_355 ? 6'h1a : _ctrlsignals_T_3680; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3682 = _ctrlsignals_T_353 ? 6'h1b : _ctrlsignals_T_3681; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3683 = _ctrlsignals_T_351 ? 6'h4 : _ctrlsignals_T_3682; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3684 = _ctrlsignals_T_349 ? 6'h6 : _ctrlsignals_T_3683; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3685 = _ctrlsignals_T_347 ? 6'h7 : _ctrlsignals_T_3684; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3686 = _ctrlsignals_T_345 ? 6'he : _ctrlsignals_T_3685; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3687 = _ctrlsignals_T_343 ? 6'he : _ctrlsignals_T_3686; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3688 = _ctrlsignals_T_341 ? 6'he : _ctrlsignals_T_3687; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3689 = _ctrlsignals_T_339 ? 6'he : _ctrlsignals_T_3688; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3690 = _ctrlsignals_T_337 ? 6'hd : _ctrlsignals_T_3689; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3691 = _ctrlsignals_T_335 ? 6'hd : _ctrlsignals_T_3690; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3692 = _ctrlsignals_T_333 ? 6'hd : _ctrlsignals_T_3691; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3693 = _ctrlsignals_T_331 ? 6'hf : _ctrlsignals_T_3692; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3694 = _ctrlsignals_T_329 ? 6'hf : _ctrlsignals_T_3693; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3695 = _ctrlsignals_T_327 ? 6'hf : _ctrlsignals_T_3694; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3696 = _ctrlsignals_T_325 ? 6'hb : _ctrlsignals_T_3695; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3697 = _ctrlsignals_T_323 ? 6'hb : _ctrlsignals_T_3696; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3698 = _ctrlsignals_T_321 ? 6'hb : _ctrlsignals_T_3697; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3699 = _ctrlsignals_T_319 ? 6'h5 : _ctrlsignals_T_3698; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3700 = _ctrlsignals_T_317 ? 6'h5 : _ctrlsignals_T_3699; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3701 = _ctrlsignals_T_315 ? 6'h5 : _ctrlsignals_T_3700; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3702 = _ctrlsignals_T_313 ? 6'h1 : _ctrlsignals_T_3701; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3703 = _ctrlsignals_T_311 ? 6'h1 : _ctrlsignals_T_3702; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3704 = _ctrlsignals_T_309 ? 6'h1 : _ctrlsignals_T_3703; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3705 = _ctrlsignals_T_307 ? 6'ha : _ctrlsignals_T_3704; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3706 = _ctrlsignals_T_305 ? 6'hb : _ctrlsignals_T_3705; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3707 = _ctrlsignals_T_303 ? 6'hb : _ctrlsignals_T_3706; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3708 = _ctrlsignals_T_301 ? 6'hb : _ctrlsignals_T_3707; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3709 = _ctrlsignals_T_299 ? 6'hc : _ctrlsignals_T_3708; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3710 = _ctrlsignals_T_297 ? 6'hc : _ctrlsignals_T_3709; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3711 = _ctrlsignals_T_295 ? 6'he : _ctrlsignals_T_3710; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3712 = _ctrlsignals_T_293 ? 6'he : _ctrlsignals_T_3711; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3713 = _ctrlsignals_T_291 ? 6'ha : _ctrlsignals_T_3712; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3714 = _ctrlsignals_T_289 ? 6'ha : _ctrlsignals_T_3713; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3715 = _ctrlsignals_T_287 ? 6'hd : _ctrlsignals_T_3714; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3716 = _ctrlsignals_T_285 ? 6'hd : _ctrlsignals_T_3715; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3717 = _ctrlsignals_T_283 ? 6'hc : _ctrlsignals_T_3716; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3718 = _ctrlsignals_T_281 ? 6'hc : _ctrlsignals_T_3717; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3719 = _ctrlsignals_T_279 ? 6'h3 : _ctrlsignals_T_3718; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3720 = _ctrlsignals_T_277 ? 6'h3 : _ctrlsignals_T_3719; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3721 = _ctrlsignals_T_275 ? 6'h3 : _ctrlsignals_T_3720; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3722 = _ctrlsignals_T_273 ? 6'h2 : _ctrlsignals_T_3721; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3723 = _ctrlsignals_T_271 ? 6'h2 : _ctrlsignals_T_3722; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3724 = _ctrlsignals_T_269 ? 6'h2 : _ctrlsignals_T_3723; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3725 = _ctrlsignals_T_267 ? 6'h4 : _ctrlsignals_T_3724; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3726 = _ctrlsignals_T_265 ? 6'h4 : _ctrlsignals_T_3725; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3727 = _ctrlsignals_T_263 ? 6'h4 : _ctrlsignals_T_3726; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3728 = _ctrlsignals_T_261 ? 6'h6 : _ctrlsignals_T_3727; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3729 = _ctrlsignals_T_259 ? 6'h6 : _ctrlsignals_T_3728; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3730 = _ctrlsignals_T_257 ? 6'h6 : _ctrlsignals_T_3729; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3731 = _ctrlsignals_T_255 ? 6'h7 : _ctrlsignals_T_3730; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3732 = _ctrlsignals_T_253 ? 6'h7 : _ctrlsignals_T_3731; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3733 = _ctrlsignals_T_251 ? 6'h7 : _ctrlsignals_T_3732; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3734 = _ctrlsignals_T_249 ? 6'h9 : _ctrlsignals_T_3733; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3735 = _ctrlsignals_T_247 ? 6'h9 : _ctrlsignals_T_3734; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3736 = _ctrlsignals_T_245 ? 6'h8 : _ctrlsignals_T_3735; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3737 = _ctrlsignals_T_243 ? 6'h8 : _ctrlsignals_T_3736; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3738 = _ctrlsignals_T_241 ? 6'ha : _ctrlsignals_T_3737; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3739 = _ctrlsignals_T_239 ? 6'ha : _ctrlsignals_T_3738; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3740 = _ctrlsignals_T_237 ? 6'ha : _ctrlsignals_T_3739; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3741 = _ctrlsignals_T_235 ? 6'ha : _ctrlsignals_T_3740; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3742 = _ctrlsignals_T_233 ? 6'h1 : _ctrlsignals_T_3741; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3743 = _ctrlsignals_T_231 ? 6'h1 : _ctrlsignals_T_3742; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3744 = _ctrlsignals_T_229 ? 6'h1 : _ctrlsignals_T_3743; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3745 = _ctrlsignals_T_227 ? 6'h0 : _ctrlsignals_T_3744; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3746 = _ctrlsignals_T_225 ? 6'h0 : _ctrlsignals_T_3745; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3747 = _ctrlsignals_T_223 ? 6'h0 : _ctrlsignals_T_3746; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3748 = _ctrlsignals_T_221 ? 6'h0 : _ctrlsignals_T_3747; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3749 = _ctrlsignals_T_219 ? 6'h0 : _ctrlsignals_T_3748; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3750 = _ctrlsignals_T_217 ? 6'h6 : _ctrlsignals_T_3749; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3751 = _ctrlsignals_T_215 ? 6'h6 : _ctrlsignals_T_3750; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3752 = _ctrlsignals_T_213 ? 6'h5 : _ctrlsignals_T_3751; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3753 = _ctrlsignals_T_211 ? 6'h5 : _ctrlsignals_T_3752; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3754 = _ctrlsignals_T_209 ? 6'h7 : _ctrlsignals_T_3753; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3755 = _ctrlsignals_T_207 ? 6'h7 : _ctrlsignals_T_3754; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3756 = _ctrlsignals_T_205 ? 6'h4 : _ctrlsignals_T_3755; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3757 = _ctrlsignals_T_203 ? 6'h4 : _ctrlsignals_T_3756; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3758 = _ctrlsignals_T_201 ? 6'h10 : _ctrlsignals_T_3757; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3759 = _ctrlsignals_T_199 ? 6'h10 : _ctrlsignals_T_3758; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3760 = _ctrlsignals_T_197 ? 6'hf : _ctrlsignals_T_3759; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3761 = _ctrlsignals_T_195 ? 6'hf : _ctrlsignals_T_3760; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3762 = _ctrlsignals_T_193 ? 6'h11 : _ctrlsignals_T_3761; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3763 = _ctrlsignals_T_191 ? 6'h11 : _ctrlsignals_T_3762; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3764 = _ctrlsignals_T_189 ? 6'he : _ctrlsignals_T_3763; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3765 = _ctrlsignals_T_187 ? 6'he : _ctrlsignals_T_3764; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3766 = _ctrlsignals_T_185 ? 6'h2 : _ctrlsignals_T_3765; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3767 = _ctrlsignals_T_183 ? 6'h2 : _ctrlsignals_T_3766; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3768 = _ctrlsignals_T_181 ? 6'h0 : _ctrlsignals_T_3767; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3769 = _ctrlsignals_T_179 ? 6'h0 : _ctrlsignals_T_3768; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3770 = _ctrlsignals_T_177 ? 6'h0 : _ctrlsignals_T_3769; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3771 = _ctrlsignals_T_175 ? 6'h0 : _ctrlsignals_T_3770; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3772 = _ctrlsignals_T_173 ? 6'h0 : _ctrlsignals_T_3771; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3773 = _ctrlsignals_T_171 ? 6'h0 : _ctrlsignals_T_3772; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3774 = _ctrlsignals_T_169 ? 6'h21 : _ctrlsignals_T_3773; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3775 = _ctrlsignals_T_167 ? 6'h20 : _ctrlsignals_T_3774; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3776 = _ctrlsignals_T_165 ? 6'h12 : _ctrlsignals_T_3775; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3777 = _ctrlsignals_T_163 ? 6'ha : _ctrlsignals_T_3776; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3778 = _ctrlsignals_T_161 ? 6'hb : _ctrlsignals_T_3777; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3779 = _ctrlsignals_T_159 ? 6'hc : _ctrlsignals_T_3778; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3780 = _ctrlsignals_T_143 ? 6'h16 : _ctrlsignals_T_3779; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3781 = _ctrlsignals_T_155 ? 6'h19 : _ctrlsignals_T_3780; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3782 = _ctrlsignals_T_153 ? 6'h18 : _ctrlsignals_T_3781; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3783 = _ctrlsignals_T_151 ? 6'h9 : _ctrlsignals_T_3782; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3784 = _ctrlsignals_T_149 ? 6'h8 : _ctrlsignals_T_3783; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3785 = _ctrlsignals_T_147 ? 6'h14 : _ctrlsignals_T_3784; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3786 = _ctrlsignals_T_145 ? 6'h15 : _ctrlsignals_T_3785; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3787 = _ctrlsignals_T_143 ? 6'h16 : _ctrlsignals_T_3786; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3788 = _ctrlsignals_T_141 ? 6'h1 : _ctrlsignals_T_3787; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3789 = _ctrlsignals_T_139 ? 6'h0 : _ctrlsignals_T_3788; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3790 = _ctrlsignals_T_137 ? 6'h2 : _ctrlsignals_T_3789; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3791 = _ctrlsignals_T_135 ? 6'h1 : _ctrlsignals_T_3790; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3792 = _ctrlsignals_T_133 ? 6'h0 : _ctrlsignals_T_3791; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3793 = _ctrlsignals_T_131 ? 6'h7 : _ctrlsignals_T_3792; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3794 = _ctrlsignals_T_129 ? 6'h6 : _ctrlsignals_T_3793; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3795 = _ctrlsignals_T_127 ? 6'h5 : _ctrlsignals_T_3794; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3796 = _ctrlsignals_T_125 ? 6'h4 : _ctrlsignals_T_3795; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3797 = _ctrlsignals_T_123 ? 6'h3 : _ctrlsignals_T_3796; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3798 = _ctrlsignals_T_121 ? 6'h1 : _ctrlsignals_T_3797; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3799 = _ctrlsignals_T_119 ? 6'h2 : _ctrlsignals_T_3798; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3800 = _ctrlsignals_T_117 ? 6'h0 : _ctrlsignals_T_3799; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3801 = _ctrlsignals_T_115 ? 6'h16 : _ctrlsignals_T_3800; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3802 = _ctrlsignals_T_113 ? 6'h17 : _ctrlsignals_T_3801; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3803 = _ctrlsignals_T_111 ? 6'h15 : _ctrlsignals_T_3802; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3804 = _ctrlsignals_T_109 ? 6'h14 : _ctrlsignals_T_3803; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3805 = _ctrlsignals_T_107 ? 6'h0 : _ctrlsignals_T_3804; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3806 = _ctrlsignals_T_105 ? 6'hb : _ctrlsignals_T_3805; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3807 = _ctrlsignals_T_103 ? 6'h5 : _ctrlsignals_T_3806; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3808 = _ctrlsignals_T_101 ? 6'h1 : _ctrlsignals_T_3807; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3809 = _ctrlsignals_T_99 ? 6'hb : _ctrlsignals_T_3808; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3810 = _ctrlsignals_T_97 ? 6'h5 : _ctrlsignals_T_3809; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3811 = _ctrlsignals_T_95 ? 6'h1 : _ctrlsignals_T_3810; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3812 = _ctrlsignals_T_93 ? 6'h4 : _ctrlsignals_T_3811; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3813 = _ctrlsignals_T_91 ? 6'h6 : _ctrlsignals_T_3812; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3814 = _ctrlsignals_T_89 ? 6'h7 : _ctrlsignals_T_3813; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3815 = _ctrlsignals_T_87 ? 6'he : _ctrlsignals_T_3814; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3816 = _ctrlsignals_T_85 ? 6'hc : _ctrlsignals_T_3815; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3817 = _ctrlsignals_T_83 ? 6'ha : _ctrlsignals_T_3816; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3818 = _ctrlsignals_T_81 ? 6'h0 : _ctrlsignals_T_3817; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3819 = _ctrlsignals_T_79 ? 6'h4 : _ctrlsignals_T_3818; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3820 = _ctrlsignals_T_77 ? 6'h6 : _ctrlsignals_T_3819; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3821 = _ctrlsignals_T_75 ? 6'h7 : _ctrlsignals_T_3820; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3822 = _ctrlsignals_T_73 ? 6'he : _ctrlsignals_T_3821; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3823 = _ctrlsignals_T_71 ? 6'hc : _ctrlsignals_T_3822; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3824 = _ctrlsignals_T_69 ? 6'h0 : _ctrlsignals_T_3823; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3825 = _ctrlsignals_T_67 ? 6'h8 : _ctrlsignals_T_3824; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3826 = _ctrlsignals_T_65 ? 6'h0 : _ctrlsignals_T_3825; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3827 = _ctrlsignals_T_63 ? 6'h0 : _ctrlsignals_T_3826; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3828 = _ctrlsignals_T_61 ? 6'h0 : _ctrlsignals_T_3827; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3829 = _ctrlsignals_T_59 ? 6'h0 : _ctrlsignals_T_3828; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3830 = _ctrlsignals_T_57 ? 6'h0 : _ctrlsignals_T_3829; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3831 = _ctrlsignals_T_55 ? 6'h0 : _ctrlsignals_T_3830; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3832 = _ctrlsignals_T_53 ? 6'h0 : _ctrlsignals_T_3831; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3833 = _ctrlsignals_T_51 ? 6'h0 : _ctrlsignals_T_3832; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3834 = _ctrlsignals_T_49 ? 6'h0 : _ctrlsignals_T_3833; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3835 = _ctrlsignals_T_47 ? 6'h0 : _ctrlsignals_T_3834; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3836 = _ctrlsignals_T_45 ? 6'h0 : _ctrlsignals_T_3835; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3837 = _ctrlsignals_T_43 ? 6'h0 : _ctrlsignals_T_3836; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3838 = _ctrlsignals_T_41 ? 6'h0 : _ctrlsignals_T_3837; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3839 = _ctrlsignals_T_39 ? 6'h0 : _ctrlsignals_T_3838; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3840 = _ctrlsignals_T_37 ? 6'h0 : _ctrlsignals_T_3839; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3841 = _ctrlsignals_T_35 ? 6'h0 : _ctrlsignals_T_3840; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3842 = _ctrlsignals_T_33 ? 6'h0 : _ctrlsignals_T_3841; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3843 = _ctrlsignals_T_31 ? 6'h0 : _ctrlsignals_T_3842; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3844 = _ctrlsignals_T_29 ? 6'hf : _ctrlsignals_T_3843; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3845 = _ctrlsignals_T_27 ? 6'hd : _ctrlsignals_T_3844; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3846 = _ctrlsignals_T_25 ? 6'he : _ctrlsignals_T_3845; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3847 = _ctrlsignals_T_23 ? 6'hc : _ctrlsignals_T_3846; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3848 = _ctrlsignals_T_21 ? 6'h2 : _ctrlsignals_T_3847; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3849 = _ctrlsignals_T_19 ? 6'h3 : _ctrlsignals_T_3848; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3850 = _ctrlsignals_T_17 ? 6'h0 : _ctrlsignals_T_3849; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3851 = _ctrlsignals_T_15 ? 6'h0 : _ctrlsignals_T_3850; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3852 = _ctrlsignals_T_13 ? 6'h0 : _ctrlsignals_T_3851; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3853 = _ctrlsignals_T_11 ? 6'hf : _ctrlsignals_T_3852; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3854 = _ctrlsignals_T_9 ? 6'hd : _ctrlsignals_T_3853; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3855 = _ctrlsignals_T_7 ? 6'he : _ctrlsignals_T_3854; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3856 = _ctrlsignals_T_5 ? 6'hc : _ctrlsignals_T_3855; // @[Lookup.scala 34:39]
  wire [5:0] _ctrlsignals_T_3857 = _ctrlsignals_T_3 ? 6'h2 : _ctrlsignals_T_3856; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4250 = _ctrlsignals_T_181 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4251 = _ctrlsignals_T_179 ? 2'h2 : _ctrlsignals_T_4250; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4252 = _ctrlsignals_T_177 ? 2'h2 : _ctrlsignals_T_4251; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4253 = _ctrlsignals_T_175 ? 2'h1 : _ctrlsignals_T_4252; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4254 = _ctrlsignals_T_173 ? 2'h1 : _ctrlsignals_T_4253; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4255 = _ctrlsignals_T_171 ? 2'h1 : _ctrlsignals_T_4254; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4256 = _ctrlsignals_T_169 ? 2'h0 : _ctrlsignals_T_4255; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4257 = _ctrlsignals_T_167 ? 2'h0 : _ctrlsignals_T_4256; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4258 = _ctrlsignals_T_165 ? 2'h0 : _ctrlsignals_T_4257; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4259 = _ctrlsignals_T_163 ? 2'h0 : _ctrlsignals_T_4258; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4260 = _ctrlsignals_T_161 ? 2'h0 : _ctrlsignals_T_4259; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4261 = _ctrlsignals_T_159 ? 2'h0 : _ctrlsignals_T_4260; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4262 = _ctrlsignals_T_143 ? 2'h0 : _ctrlsignals_T_4261; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4263 = _ctrlsignals_T_155 ? 2'h0 : _ctrlsignals_T_4262; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4264 = _ctrlsignals_T_153 ? 2'h0 : _ctrlsignals_T_4263; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4265 = _ctrlsignals_T_151 ? 2'h0 : _ctrlsignals_T_4264; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4266 = _ctrlsignals_T_149 ? 2'h0 : _ctrlsignals_T_4265; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4267 = _ctrlsignals_T_147 ? 2'h0 : _ctrlsignals_T_4266; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4268 = _ctrlsignals_T_145 ? 2'h0 : _ctrlsignals_T_4267; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4269 = _ctrlsignals_T_143 ? 2'h0 : _ctrlsignals_T_4268; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4270 = _ctrlsignals_T_141 ? 2'h0 : _ctrlsignals_T_4269; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4271 = _ctrlsignals_T_139 ? 2'h0 : _ctrlsignals_T_4270; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4272 = _ctrlsignals_T_137 ? 2'h0 : _ctrlsignals_T_4271; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4273 = _ctrlsignals_T_135 ? 2'h0 : _ctrlsignals_T_4272; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4274 = _ctrlsignals_T_133 ? 2'h0 : _ctrlsignals_T_4273; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4275 = _ctrlsignals_T_131 ? 2'h0 : _ctrlsignals_T_4274; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4276 = _ctrlsignals_T_129 ? 2'h0 : _ctrlsignals_T_4275; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4277 = _ctrlsignals_T_127 ? 2'h0 : _ctrlsignals_T_4276; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4278 = _ctrlsignals_T_125 ? 2'h0 : _ctrlsignals_T_4277; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4279 = _ctrlsignals_T_123 ? 2'h0 : _ctrlsignals_T_4278; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4280 = _ctrlsignals_T_121 ? 2'h0 : _ctrlsignals_T_4279; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4281 = _ctrlsignals_T_119 ? 2'h0 : _ctrlsignals_T_4280; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4282 = _ctrlsignals_T_117 ? 2'h0 : _ctrlsignals_T_4281; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4283 = _ctrlsignals_T_115 ? 2'h0 : _ctrlsignals_T_4282; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4284 = _ctrlsignals_T_113 ? 2'h0 : _ctrlsignals_T_4283; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4285 = _ctrlsignals_T_111 ? 2'h0 : _ctrlsignals_T_4284; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4286 = _ctrlsignals_T_109 ? 2'h0 : _ctrlsignals_T_4285; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4287 = _ctrlsignals_T_107 ? 2'h0 : _ctrlsignals_T_4286; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4288 = _ctrlsignals_T_105 ? 2'h0 : _ctrlsignals_T_4287; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4289 = _ctrlsignals_T_103 ? 2'h0 : _ctrlsignals_T_4288; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4290 = _ctrlsignals_T_101 ? 2'h0 : _ctrlsignals_T_4289; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4291 = _ctrlsignals_T_99 ? 2'h0 : _ctrlsignals_T_4290; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4292 = _ctrlsignals_T_97 ? 2'h0 : _ctrlsignals_T_4291; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4293 = _ctrlsignals_T_95 ? 2'h0 : _ctrlsignals_T_4292; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4294 = _ctrlsignals_T_93 ? 2'h0 : _ctrlsignals_T_4293; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4295 = _ctrlsignals_T_91 ? 2'h0 : _ctrlsignals_T_4294; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4296 = _ctrlsignals_T_89 ? 2'h0 : _ctrlsignals_T_4295; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4297 = _ctrlsignals_T_87 ? 2'h0 : _ctrlsignals_T_4296; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4298 = _ctrlsignals_T_85 ? 2'h0 : _ctrlsignals_T_4297; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4299 = _ctrlsignals_T_83 ? 2'h0 : _ctrlsignals_T_4298; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4300 = _ctrlsignals_T_81 ? 2'h0 : _ctrlsignals_T_4299; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4301 = _ctrlsignals_T_79 ? 2'h0 : _ctrlsignals_T_4300; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4302 = _ctrlsignals_T_77 ? 2'h0 : _ctrlsignals_T_4301; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4303 = _ctrlsignals_T_75 ? 2'h0 : _ctrlsignals_T_4302; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4304 = _ctrlsignals_T_73 ? 2'h0 : _ctrlsignals_T_4303; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4305 = _ctrlsignals_T_71 ? 2'h0 : _ctrlsignals_T_4304; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4306 = _ctrlsignals_T_69 ? 2'h0 : _ctrlsignals_T_4305; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4307 = _ctrlsignals_T_67 ? 2'h0 : _ctrlsignals_T_4306; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4308 = _ctrlsignals_T_65 ? 2'h2 : _ctrlsignals_T_4307; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4309 = _ctrlsignals_T_63 ? 2'h2 : _ctrlsignals_T_4308; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4310 = _ctrlsignals_T_61 ? 2'h2 : _ctrlsignals_T_4309; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4311 = _ctrlsignals_T_59 ? 2'h1 : _ctrlsignals_T_4310; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4312 = _ctrlsignals_T_57 ? 2'h1 : _ctrlsignals_T_4311; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4313 = _ctrlsignals_T_55 ? 2'h1 : _ctrlsignals_T_4312; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4314 = _ctrlsignals_T_53 ? 2'h1 : _ctrlsignals_T_4313; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4315 = _ctrlsignals_T_51 ? 2'h1 : _ctrlsignals_T_4314; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4316 = _ctrlsignals_T_49 ? 2'h0 : _ctrlsignals_T_4315; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4317 = _ctrlsignals_T_47 ? 2'h0 : _ctrlsignals_T_4316; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4318 = _ctrlsignals_T_45 ? 2'h0 : _ctrlsignals_T_4317; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4319 = _ctrlsignals_T_43 ? 2'h0 : _ctrlsignals_T_4318; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4320 = _ctrlsignals_T_41 ? 2'h0 : _ctrlsignals_T_4319; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4321 = _ctrlsignals_T_39 ? 2'h0 : _ctrlsignals_T_4320; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4322 = _ctrlsignals_T_37 ? 2'h0 : _ctrlsignals_T_4321; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4323 = _ctrlsignals_T_35 ? 2'h0 : _ctrlsignals_T_4322; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4324 = _ctrlsignals_T_33 ? 2'h0 : _ctrlsignals_T_4323; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4325 = _ctrlsignals_T_31 ? 2'h0 : _ctrlsignals_T_4324; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4326 = _ctrlsignals_T_29 ? 2'h0 : _ctrlsignals_T_4325; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4327 = _ctrlsignals_T_27 ? 2'h0 : _ctrlsignals_T_4326; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4328 = _ctrlsignals_T_25 ? 2'h0 : _ctrlsignals_T_4327; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4329 = _ctrlsignals_T_23 ? 2'h0 : _ctrlsignals_T_4328; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4330 = _ctrlsignals_T_21 ? 2'h0 : _ctrlsignals_T_4329; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4331 = _ctrlsignals_T_19 ? 2'h0 : _ctrlsignals_T_4330; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4332 = _ctrlsignals_T_17 ? 2'h0 : _ctrlsignals_T_4331; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4333 = _ctrlsignals_T_15 ? 2'h0 : _ctrlsignals_T_4332; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4334 = _ctrlsignals_T_13 ? 2'h0 : _ctrlsignals_T_4333; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4335 = _ctrlsignals_T_11 ? 2'h0 : _ctrlsignals_T_4334; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4336 = _ctrlsignals_T_9 ? 2'h0 : _ctrlsignals_T_4335; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4337 = _ctrlsignals_T_7 ? 2'h0 : _ctrlsignals_T_4336; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4338 = _ctrlsignals_T_5 ? 2'h0 : _ctrlsignals_T_4337; // @[Lookup.scala 34:39]
  wire [1:0] _ctrlsignals_T_4339 = _ctrlsignals_T_3 ? 2'h0 : _ctrlsignals_T_4338; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4554 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_57 | _ctrlsignals_T_59; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4555 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_4554; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4556 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_4555; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4557 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_4556; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4558 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_4557; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4559 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_4558; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4560 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_4559; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4561 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_4560; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4562 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_4561; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4563 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_4562; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4564 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_4563; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4565 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_4564; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4566 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_4565; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4567 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_4566; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4568 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_4567; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4569 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_4568; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4570 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_4569; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4571 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_4570; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4572 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_4571; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4573 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_4572; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4574 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_4573; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4575 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_4574; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4576 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_4575; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4577 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_4576; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4578 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_4577; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4579 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_4578; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4580 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_4579; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4799 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_49; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4800 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_4799; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4801 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_4800; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4802 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_4801; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4803 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_4802; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4804 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_4803; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4805 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_4804; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4806 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_4805; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4807 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_4806; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4808 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_4807; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4809 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_4808; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4810 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_4809; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4811 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_4810; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4812 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_4811; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4813 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_4812; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4814 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_4813; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4815 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_4814; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4816 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_4815; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4817 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_4816; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4818 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_4817; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4819 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_4818; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4820 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_4819; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4821 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_4820; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4863 = _ctrlsignals_T_401 ? 1'h0 : _ctrlsignals_T_403 | (_ctrlsignals_T_405 | (_ctrlsignals_T_407
     | (_ctrlsignals_T_409 | (_ctrlsignals_T_411 | (_ctrlsignals_T_413 | (_ctrlsignals_T_415 | (_ctrlsignals_T_417 | (
    _ctrlsignals_T_419 | (_ctrlsignals_T_421 | (_ctrlsignals_T_423 | _ctrlsignals_T_425)))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4864 = _ctrlsignals_T_399 ? 1'h0 : _ctrlsignals_T_4863; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4865 = _ctrlsignals_T_397 ? 1'h0 : _ctrlsignals_T_4864; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4866 = _ctrlsignals_T_395 ? 1'h0 : _ctrlsignals_T_4865; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4867 = _ctrlsignals_T_393 ? 1'h0 : _ctrlsignals_T_4866; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4868 = _ctrlsignals_T_391 ? 1'h0 : _ctrlsignals_T_4867; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4869 = _ctrlsignals_T_389 ? 1'h0 : _ctrlsignals_T_4868; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4870 = _ctrlsignals_T_387 ? 1'h0 : _ctrlsignals_T_4869; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4871 = _ctrlsignals_T_385 ? 1'h0 : _ctrlsignals_T_4870; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4872 = _ctrlsignals_T_383 ? 1'h0 : _ctrlsignals_T_4871; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4873 = _ctrlsignals_T_381 ? 1'h0 : _ctrlsignals_T_4872; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4874 = _ctrlsignals_T_379 ? 1'h0 : _ctrlsignals_T_4873; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4875 = _ctrlsignals_T_377 ? 1'h0 : _ctrlsignals_T_4874; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4876 = _ctrlsignals_T_375 ? 1'h0 : _ctrlsignals_T_4875; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4877 = _ctrlsignals_T_373 ? 1'h0 : _ctrlsignals_T_4876; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4878 = _ctrlsignals_T_371 ? 1'h0 : _ctrlsignals_T_4877; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4879 = _ctrlsignals_T_369 ? 1'h0 : _ctrlsignals_T_4878; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4880 = _ctrlsignals_T_367 ? 1'h0 : _ctrlsignals_T_4879; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4881 = _ctrlsignals_T_365 ? 1'h0 : _ctrlsignals_T_4880; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4882 = _ctrlsignals_T_363 ? 1'h0 : _ctrlsignals_T_4881; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4883 = _ctrlsignals_T_361 ? 1'h0 : _ctrlsignals_T_4882; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4884 = _ctrlsignals_T_359 ? 1'h0 : _ctrlsignals_T_4883; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4885 = _ctrlsignals_T_357 ? 1'h0 : _ctrlsignals_T_4884; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4886 = _ctrlsignals_T_355 ? 1'h0 : _ctrlsignals_T_4885; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4887 = _ctrlsignals_T_353 ? 1'h0 : _ctrlsignals_T_4886; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4888 = _ctrlsignals_T_351 ? 1'h0 : _ctrlsignals_T_4887; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4889 = _ctrlsignals_T_349 ? 1'h0 : _ctrlsignals_T_4888; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4890 = _ctrlsignals_T_347 ? 1'h0 : _ctrlsignals_T_4889; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4891 = _ctrlsignals_T_345 ? 1'h0 : _ctrlsignals_T_4890; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4892 = _ctrlsignals_T_343 ? 1'h0 : _ctrlsignals_T_4891; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4893 = _ctrlsignals_T_341 ? 1'h0 : _ctrlsignals_T_4892; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4894 = _ctrlsignals_T_339 ? 1'h0 : _ctrlsignals_T_4893; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4895 = _ctrlsignals_T_337 ? 1'h0 : _ctrlsignals_T_4894; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4896 = _ctrlsignals_T_335 ? 1'h0 : _ctrlsignals_T_4895; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4897 = _ctrlsignals_T_333 ? 1'h0 : _ctrlsignals_T_4896; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4898 = _ctrlsignals_T_331 ? 1'h0 : _ctrlsignals_T_4897; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4899 = _ctrlsignals_T_329 ? 1'h0 : _ctrlsignals_T_4898; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4900 = _ctrlsignals_T_327 ? 1'h0 : _ctrlsignals_T_4899; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4901 = _ctrlsignals_T_325 ? 1'h0 : _ctrlsignals_T_4900; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4902 = _ctrlsignals_T_323 ? 1'h0 : _ctrlsignals_T_4901; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4903 = _ctrlsignals_T_321 ? 1'h0 : _ctrlsignals_T_4902; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4904 = _ctrlsignals_T_319 ? 1'h0 : _ctrlsignals_T_4903; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4905 = _ctrlsignals_T_317 ? 1'h0 : _ctrlsignals_T_4904; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4906 = _ctrlsignals_T_315 ? 1'h0 : _ctrlsignals_T_4905; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4907 = _ctrlsignals_T_313 ? 1'h0 : _ctrlsignals_T_4906; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4908 = _ctrlsignals_T_311 ? 1'h0 : _ctrlsignals_T_4907; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4909 = _ctrlsignals_T_309 ? 1'h0 : _ctrlsignals_T_4908; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4910 = _ctrlsignals_T_307 ? 1'h0 : _ctrlsignals_T_4909; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4911 = _ctrlsignals_T_305 ? 1'h0 : _ctrlsignals_T_4910; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4912 = _ctrlsignals_T_303 ? 1'h0 : _ctrlsignals_T_4911; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4913 = _ctrlsignals_T_301 ? 1'h0 : _ctrlsignals_T_4912; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4914 = _ctrlsignals_T_299 ? 1'h0 : _ctrlsignals_T_4913; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4915 = _ctrlsignals_T_297 ? 1'h0 : _ctrlsignals_T_4914; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4916 = _ctrlsignals_T_295 ? 1'h0 : _ctrlsignals_T_4915; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4917 = _ctrlsignals_T_293 ? 1'h0 : _ctrlsignals_T_4916; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4918 = _ctrlsignals_T_291 ? 1'h0 : _ctrlsignals_T_4917; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4919 = _ctrlsignals_T_289 ? 1'h0 : _ctrlsignals_T_4918; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4920 = _ctrlsignals_T_287 ? 1'h0 : _ctrlsignals_T_4919; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4921 = _ctrlsignals_T_285 ? 1'h0 : _ctrlsignals_T_4920; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4922 = _ctrlsignals_T_283 ? 1'h0 : _ctrlsignals_T_4921; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4923 = _ctrlsignals_T_281 ? 1'h0 : _ctrlsignals_T_4922; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4924 = _ctrlsignals_T_279 ? 1'h0 : _ctrlsignals_T_4923; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4925 = _ctrlsignals_T_277 ? 1'h0 : _ctrlsignals_T_4924; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4926 = _ctrlsignals_T_275 ? 1'h0 : _ctrlsignals_T_4925; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4927 = _ctrlsignals_T_273 ? 1'h0 : _ctrlsignals_T_4926; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4928 = _ctrlsignals_T_271 ? 1'h0 : _ctrlsignals_T_4927; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4929 = _ctrlsignals_T_269 ? 1'h0 : _ctrlsignals_T_4928; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4930 = _ctrlsignals_T_267 ? 1'h0 : _ctrlsignals_T_4929; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4931 = _ctrlsignals_T_265 ? 1'h0 : _ctrlsignals_T_4930; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4932 = _ctrlsignals_T_263 ? 1'h0 : _ctrlsignals_T_4931; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4933 = _ctrlsignals_T_261 ? 1'h0 : _ctrlsignals_T_4932; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4934 = _ctrlsignals_T_259 ? 1'h0 : _ctrlsignals_T_4933; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4935 = _ctrlsignals_T_257 ? 1'h0 : _ctrlsignals_T_4934; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4936 = _ctrlsignals_T_255 ? 1'h0 : _ctrlsignals_T_4935; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4937 = _ctrlsignals_T_253 ? 1'h0 : _ctrlsignals_T_4936; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4938 = _ctrlsignals_T_251 ? 1'h0 : _ctrlsignals_T_4937; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4939 = _ctrlsignals_T_249 ? 1'h0 : _ctrlsignals_T_4938; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4940 = _ctrlsignals_T_247 ? 1'h0 : _ctrlsignals_T_4939; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4941 = _ctrlsignals_T_245 ? 1'h0 : _ctrlsignals_T_4940; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4942 = _ctrlsignals_T_243 ? 1'h0 : _ctrlsignals_T_4941; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4943 = _ctrlsignals_T_241 ? 1'h0 : _ctrlsignals_T_4942; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4944 = _ctrlsignals_T_239 ? 1'h0 : _ctrlsignals_T_4943; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4945 = _ctrlsignals_T_237 ? 1'h0 : _ctrlsignals_T_4944; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4946 = _ctrlsignals_T_235 ? 1'h0 : _ctrlsignals_T_4945; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4947 = _ctrlsignals_T_233 ? 1'h0 : _ctrlsignals_T_4946; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4948 = _ctrlsignals_T_231 ? 1'h0 : _ctrlsignals_T_4947; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4949 = _ctrlsignals_T_229 ? 1'h0 : _ctrlsignals_T_4948; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4950 = _ctrlsignals_T_227 ? 1'h0 : _ctrlsignals_T_4949; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4951 = _ctrlsignals_T_225 ? 1'h0 : _ctrlsignals_T_4950; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4952 = _ctrlsignals_T_223 ? 1'h0 : _ctrlsignals_T_4951; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4953 = _ctrlsignals_T_221 ? 1'h0 : _ctrlsignals_T_4952; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4954 = _ctrlsignals_T_219 ? 1'h0 : _ctrlsignals_T_4953; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4955 = _ctrlsignals_T_217 ? 1'h0 : _ctrlsignals_T_4954; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4956 = _ctrlsignals_T_215 ? 1'h0 : _ctrlsignals_T_4955; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4957 = _ctrlsignals_T_213 ? 1'h0 : _ctrlsignals_T_4956; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4958 = _ctrlsignals_T_211 ? 1'h0 : _ctrlsignals_T_4957; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4959 = _ctrlsignals_T_209 ? 1'h0 : _ctrlsignals_T_4958; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4960 = _ctrlsignals_T_207 ? 1'h0 : _ctrlsignals_T_4959; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4961 = _ctrlsignals_T_205 ? 1'h0 : _ctrlsignals_T_4960; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4962 = _ctrlsignals_T_203 ? 1'h0 : _ctrlsignals_T_4961; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4963 = _ctrlsignals_T_201 ? 1'h0 : _ctrlsignals_T_4962; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4964 = _ctrlsignals_T_199 ? 1'h0 : _ctrlsignals_T_4963; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4965 = _ctrlsignals_T_197 ? 1'h0 : _ctrlsignals_T_4964; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4966 = _ctrlsignals_T_195 ? 1'h0 : _ctrlsignals_T_4965; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4967 = _ctrlsignals_T_193 ? 1'h0 : _ctrlsignals_T_4966; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4968 = _ctrlsignals_T_191 ? 1'h0 : _ctrlsignals_T_4967; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4969 = _ctrlsignals_T_189 ? 1'h0 : _ctrlsignals_T_4968; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4970 = _ctrlsignals_T_187 ? 1'h0 : _ctrlsignals_T_4969; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4971 = _ctrlsignals_T_185 ? 1'h0 : _ctrlsignals_T_4970; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4972 = _ctrlsignals_T_183 ? 1'h0 : _ctrlsignals_T_4971; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4973 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_4972; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4974 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_4973; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4975 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_4974; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4976 = _ctrlsignals_T_175 ? 1'h0 : _ctrlsignals_T_4975; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4977 = _ctrlsignals_T_173 ? 1'h0 : _ctrlsignals_T_4976; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4978 = _ctrlsignals_T_171 ? 1'h0 : _ctrlsignals_T_4977; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4979 = _ctrlsignals_T_169 ? 1'h0 : _ctrlsignals_T_4978; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4980 = _ctrlsignals_T_167 ? 1'h0 : _ctrlsignals_T_4979; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4981 = _ctrlsignals_T_165 ? 1'h0 : _ctrlsignals_T_4980; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4982 = _ctrlsignals_T_163 ? 1'h0 : _ctrlsignals_T_4981; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4983 = _ctrlsignals_T_161 ? 1'h0 : _ctrlsignals_T_4982; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4984 = _ctrlsignals_T_159 ? 1'h0 : _ctrlsignals_T_4983; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4985 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_4984; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4986 = _ctrlsignals_T_155 ? 1'h0 : _ctrlsignals_T_4985; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4987 = _ctrlsignals_T_153 ? 1'h0 : _ctrlsignals_T_4986; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4988 = _ctrlsignals_T_151 ? 1'h0 : _ctrlsignals_T_4987; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4989 = _ctrlsignals_T_149 ? 1'h0 : _ctrlsignals_T_4988; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4990 = _ctrlsignals_T_147 ? 1'h0 : _ctrlsignals_T_4989; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4991 = _ctrlsignals_T_145 ? 1'h0 : _ctrlsignals_T_4990; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4992 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_4991; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4995 = _ctrlsignals_T_137 ? 1'h0 : _ctrlsignals_T_139 | (_ctrlsignals_T_141 | _ctrlsignals_T_4992
    ); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4996 = _ctrlsignals_T_135 ? 1'h0 : _ctrlsignals_T_4995; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4997 = _ctrlsignals_T_133 ? 1'h0 : _ctrlsignals_T_4996; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4998 = _ctrlsignals_T_131 ? 1'h0 : _ctrlsignals_T_4997; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_4999 = _ctrlsignals_T_129 ? 1'h0 : _ctrlsignals_T_4998; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5000 = _ctrlsignals_T_127 ? 1'h0 : _ctrlsignals_T_4999; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5001 = _ctrlsignals_T_125 ? 1'h0 : _ctrlsignals_T_5000; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5006 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_117 | (_ctrlsignals_T_119 | (_ctrlsignals_T_121
     | (_ctrlsignals_T_123 | _ctrlsignals_T_5001))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5007 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_5006; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5008 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_5007; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5009 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_5008; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5010 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_5009; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5011 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_5010; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5012 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_5011; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5013 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_5012; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5014 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_5013; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5015 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_5014; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5016 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_5015; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5017 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_5016; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5018 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_5017; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5019 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_5018; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5020 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_5019; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5021 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_5020; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5022 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_5021; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5023 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_5022; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5024 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_5023; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5025 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_5024; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5026 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_5025; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5027 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_5026; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5028 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_5027; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5029 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_5028; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5030 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_5029; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5031 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_5030; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5032 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_5031; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5033 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_5032; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5034 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_5033; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5035 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_5034; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5036 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_5035; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5037 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_5036; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5038 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_5037; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5039 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_5038; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5040 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_5039; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5041 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_5040; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5042 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_5041; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5043 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_5042; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5044 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_5043; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5045 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_5044; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5046 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_5045; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5047 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_5046; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5048 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_5047; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5049 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_5048; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5050 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_5049; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5051 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_5050; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5052 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_5051; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5053 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_5052; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5054 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_5053; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5055 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_5054; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5056 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_5055; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5057 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_5056; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5058 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_5057; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5059 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_5058; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5060 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_5059; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5061 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_5060; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5062 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_5061; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5097 = _ctrlsignals_T_415 | (_ctrlsignals_T_417 | (_ctrlsignals_T_419 | (_ctrlsignals_T_421 | (
    _ctrlsignals_T_423 | (_ctrlsignals_T_425 | (_ctrlsignals_T_427 | (_ctrlsignals_T_429 | (_ctrlsignals_T_431 | (
    _ctrlsignals_T_433 | (_ctrlsignals_T_435 | (_ctrlsignals_T_437 | (_ctrlsignals_T_439 | (_ctrlsignals_T_441 | (
    _ctrlsignals_T_443 | (_ctrlsignals_T_445 | (_ctrlsignals_T_447 | (_ctrlsignals_T_449 | (_ctrlsignals_T_451 | (
    _ctrlsignals_T_453 | (_ctrlsignals_T_443 | (_ctrlsignals_T_445 | (_ctrlsignals_T_459 | (_ctrlsignals_T_461 | (
    _ctrlsignals_T_463 | (_ctrlsignals_T_465 | (_ctrlsignals_T_467 | (_ctrlsignals_T_469 | (_ctrlsignals_T_471 | (
    _ctrlsignals_T_473 | _ctrlsignals_T_475))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5127 = _ctrlsignals_T_355 | (_ctrlsignals_T_357 | (_ctrlsignals_T_359 | (_ctrlsignals_T_361 | (
    _ctrlsignals_T_363 | (_ctrlsignals_T_365 | (_ctrlsignals_T_367 | (_ctrlsignals_T_369 | (_ctrlsignals_T_371 | (
    _ctrlsignals_T_373 | (_ctrlsignals_T_375 | (_ctrlsignals_T_377 | (_ctrlsignals_T_379 | (_ctrlsignals_T_381 | (
    _ctrlsignals_T_383 | (_ctrlsignals_T_385 | (_ctrlsignals_T_387 | (_ctrlsignals_T_389 | (_ctrlsignals_T_391 | (
    _ctrlsignals_T_393 | (_ctrlsignals_T_395 | (_ctrlsignals_T_397 | (_ctrlsignals_T_399 | (_ctrlsignals_T_401 | (
    _ctrlsignals_T_403 | (_ctrlsignals_T_405 | (_ctrlsignals_T_407 | (_ctrlsignals_T_409 | (_ctrlsignals_T_411 | (
    _ctrlsignals_T_413 | _ctrlsignals_T_5097))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5157 = _ctrlsignals_T_295 | (_ctrlsignals_T_297 | (_ctrlsignals_T_299 | (_ctrlsignals_T_301 | (
    _ctrlsignals_T_303 | (_ctrlsignals_T_305 | (_ctrlsignals_T_307 | (_ctrlsignals_T_309 | (_ctrlsignals_T_311 | (
    _ctrlsignals_T_313 | (_ctrlsignals_T_315 | (_ctrlsignals_T_317 | (_ctrlsignals_T_319 | (_ctrlsignals_T_321 | (
    _ctrlsignals_T_323 | (_ctrlsignals_T_325 | (_ctrlsignals_T_327 | (_ctrlsignals_T_329 | (_ctrlsignals_T_331 | (
    _ctrlsignals_T_333 | (_ctrlsignals_T_335 | (_ctrlsignals_T_337 | (_ctrlsignals_T_339 | (_ctrlsignals_T_341 | (
    _ctrlsignals_T_343 | (_ctrlsignals_T_345 | (_ctrlsignals_T_347 | (_ctrlsignals_T_349 | (_ctrlsignals_T_351 | (
    _ctrlsignals_T_353 | _ctrlsignals_T_5127))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5187 = _ctrlsignals_T_235 | (_ctrlsignals_T_237 | (_ctrlsignals_T_239 | (_ctrlsignals_T_241 | (
    _ctrlsignals_T_243 | (_ctrlsignals_T_245 | (_ctrlsignals_T_247 | (_ctrlsignals_T_249 | (_ctrlsignals_T_251 | (
    _ctrlsignals_T_253 | (_ctrlsignals_T_255 | (_ctrlsignals_T_257 | (_ctrlsignals_T_259 | (_ctrlsignals_T_261 | (
    _ctrlsignals_T_263 | (_ctrlsignals_T_265 | (_ctrlsignals_T_267 | (_ctrlsignals_T_269 | (_ctrlsignals_T_271 | (
    _ctrlsignals_T_273 | (_ctrlsignals_T_275 | (_ctrlsignals_T_277 | (_ctrlsignals_T_279 | (_ctrlsignals_T_281 | (
    _ctrlsignals_T_283 | (_ctrlsignals_T_285 | (_ctrlsignals_T_287 | (_ctrlsignals_T_289 | (_ctrlsignals_T_291 | (
    _ctrlsignals_T_293 | _ctrlsignals_T_5157))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5214 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_183 | (_ctrlsignals_T_185 | (_ctrlsignals_T_187
     | (_ctrlsignals_T_189 | (_ctrlsignals_T_191 | (_ctrlsignals_T_193 | (_ctrlsignals_T_195 | (_ctrlsignals_T_197 | (
    _ctrlsignals_T_199 | (_ctrlsignals_T_201 | (_ctrlsignals_T_203 | (_ctrlsignals_T_205 | (_ctrlsignals_T_207 | (
    _ctrlsignals_T_209 | (_ctrlsignals_T_211 | (_ctrlsignals_T_213 | (_ctrlsignals_T_215 | (_ctrlsignals_T_217 | (
    _ctrlsignals_T_219 | (_ctrlsignals_T_221 | (_ctrlsignals_T_223 | (_ctrlsignals_T_225 | (_ctrlsignals_T_227 | (
    _ctrlsignals_T_229 | (_ctrlsignals_T_231 | (_ctrlsignals_T_233 | _ctrlsignals_T_5187))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5215 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_5214; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5216 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_5215; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5220 = _ctrlsignals_T_169 ? 1'h0 : _ctrlsignals_T_171 | (_ctrlsignals_T_173 | (_ctrlsignals_T_175
     | _ctrlsignals_T_5216)); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5221 = _ctrlsignals_T_167 ? 1'h0 : _ctrlsignals_T_5220; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5222 = _ctrlsignals_T_165 ? 1'h0 : _ctrlsignals_T_5221; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5223 = _ctrlsignals_T_163 ? 1'h0 : _ctrlsignals_T_5222; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5224 = _ctrlsignals_T_161 ? 1'h0 : _ctrlsignals_T_5223; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5225 = _ctrlsignals_T_159 ? 1'h0 : _ctrlsignals_T_5224; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5226 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_5225; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5227 = _ctrlsignals_T_155 ? 1'h0 : _ctrlsignals_T_5226; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5228 = _ctrlsignals_T_153 ? 1'h0 : _ctrlsignals_T_5227; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5229 = _ctrlsignals_T_151 ? 1'h0 : _ctrlsignals_T_5228; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5230 = _ctrlsignals_T_149 ? 1'h0 : _ctrlsignals_T_5229; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5231 = _ctrlsignals_T_147 ? 1'h0 : _ctrlsignals_T_5230; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5232 = _ctrlsignals_T_145 ? 1'h0 : _ctrlsignals_T_5231; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5233 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_5232; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5234 = _ctrlsignals_T_141 ? 1'h0 : _ctrlsignals_T_5233; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5235 = _ctrlsignals_T_139 ? 1'h0 : _ctrlsignals_T_5234; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5236 = _ctrlsignals_T_137 ? 1'h0 : _ctrlsignals_T_5235; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5237 = _ctrlsignals_T_135 ? 1'h0 : _ctrlsignals_T_5236; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5238 = _ctrlsignals_T_133 ? 1'h0 : _ctrlsignals_T_5237; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5239 = _ctrlsignals_T_131 ? 1'h0 : _ctrlsignals_T_5238; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5240 = _ctrlsignals_T_129 ? 1'h0 : _ctrlsignals_T_5239; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5241 = _ctrlsignals_T_127 ? 1'h0 : _ctrlsignals_T_5240; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5242 = _ctrlsignals_T_125 ? 1'h0 : _ctrlsignals_T_5241; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5243 = _ctrlsignals_T_123 ? 1'h0 : _ctrlsignals_T_5242; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5244 = _ctrlsignals_T_121 ? 1'h0 : _ctrlsignals_T_5243; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5245 = _ctrlsignals_T_119 ? 1'h0 : _ctrlsignals_T_5244; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5246 = _ctrlsignals_T_117 ? 1'h0 : _ctrlsignals_T_5245; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5247 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_5246; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5248 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_5247; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5249 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_5248; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5250 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_5249; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5251 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_5250; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5252 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_5251; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5253 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_5252; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5254 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_5253; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5255 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_5254; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5256 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_5255; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5257 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_5256; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5258 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_5257; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5259 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_5258; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5260 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_5259; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5261 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_5260; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5262 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_5261; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5263 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_5262; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5264 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_5263; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5265 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_5264; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5266 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_5265; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5267 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_5266; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5268 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_5267; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5269 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_5268; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5270 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_5269; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5271 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_5270; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5272 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_5271; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5273 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_5272; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5274 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_5273; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5275 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_5274; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5276 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_5275; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5277 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_5276; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5278 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_5277; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5279 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_5278; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5280 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_5279; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5281 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_5280; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5282 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_5281; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5283 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_5282; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5284 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_5283; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5285 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_5284; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5286 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_5285; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5287 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_5286; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5288 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_5287; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5289 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_5288; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5290 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_5289; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5291 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_5290; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5292 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_5291; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5293 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_5292; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5294 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_5293; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5295 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_5294; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5296 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_5295; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5297 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_5296; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5298 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_5297; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5299 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_5298; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5300 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_5299; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5301 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_5300; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5302 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_5301; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5303 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_5302; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5373 = _ctrlsignals_T_345 ? 1'h0 : _ctrlsignals_T_347 | (_ctrlsignals_T_349 | (_ctrlsignals_T_351
     | (_ctrlsignals_T_353 | (_ctrlsignals_T_355 | (_ctrlsignals_T_357 | (_ctrlsignals_T_359 | _ctrlsignals_T_361)))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5374 = _ctrlsignals_T_343 ? 1'h0 : _ctrlsignals_T_5373; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5375 = _ctrlsignals_T_341 ? 1'h0 : _ctrlsignals_T_5374; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5376 = _ctrlsignals_T_339 ? 1'h0 : _ctrlsignals_T_5375; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5377 = _ctrlsignals_T_337 ? 1'h0 : _ctrlsignals_T_5376; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5378 = _ctrlsignals_T_335 ? 1'h0 : _ctrlsignals_T_5377; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5379 = _ctrlsignals_T_333 ? 1'h0 : _ctrlsignals_T_5378; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5380 = _ctrlsignals_T_331 ? 1'h0 : _ctrlsignals_T_5379; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5381 = _ctrlsignals_T_329 ? 1'h0 : _ctrlsignals_T_5380; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5382 = _ctrlsignals_T_327 ? 1'h0 : _ctrlsignals_T_5381; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5383 = _ctrlsignals_T_325 ? 1'h0 : _ctrlsignals_T_5382; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5384 = _ctrlsignals_T_323 ? 1'h0 : _ctrlsignals_T_5383; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5385 = _ctrlsignals_T_321 ? 1'h0 : _ctrlsignals_T_5384; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5386 = _ctrlsignals_T_319 ? 1'h0 : _ctrlsignals_T_5385; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5387 = _ctrlsignals_T_317 ? 1'h0 : _ctrlsignals_T_5386; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5388 = _ctrlsignals_T_315 ? 1'h0 : _ctrlsignals_T_5387; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5389 = _ctrlsignals_T_313 ? 1'h0 : _ctrlsignals_T_5388; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5390 = _ctrlsignals_T_311 ? 1'h0 : _ctrlsignals_T_5389; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5391 = _ctrlsignals_T_309 ? 1'h0 : _ctrlsignals_T_5390; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5392 = _ctrlsignals_T_307 ? 1'h0 : _ctrlsignals_T_5391; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5393 = _ctrlsignals_T_305 ? 1'h0 : _ctrlsignals_T_5392; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5394 = _ctrlsignals_T_303 ? 1'h0 : _ctrlsignals_T_5393; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5395 = _ctrlsignals_T_301 ? 1'h0 : _ctrlsignals_T_5394; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5396 = _ctrlsignals_T_299 ? 1'h0 : _ctrlsignals_T_5395; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5397 = _ctrlsignals_T_297 ? 1'h0 : _ctrlsignals_T_5396; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5398 = _ctrlsignals_T_295 ? 1'h0 : _ctrlsignals_T_5397; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5399 = _ctrlsignals_T_293 ? 1'h0 : _ctrlsignals_T_5398; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5400 = _ctrlsignals_T_291 ? 1'h0 : _ctrlsignals_T_5399; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5401 = _ctrlsignals_T_289 ? 1'h0 : _ctrlsignals_T_5400; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5402 = _ctrlsignals_T_287 ? 1'h0 : _ctrlsignals_T_5401; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5403 = _ctrlsignals_T_285 ? 1'h0 : _ctrlsignals_T_5402; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5404 = _ctrlsignals_T_283 ? 1'h0 : _ctrlsignals_T_5403; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5405 = _ctrlsignals_T_281 ? 1'h0 : _ctrlsignals_T_5404; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5406 = _ctrlsignals_T_279 ? 1'h0 : _ctrlsignals_T_5405; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5407 = _ctrlsignals_T_277 ? 1'h0 : _ctrlsignals_T_5406; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5408 = _ctrlsignals_T_275 ? 1'h0 : _ctrlsignals_T_5407; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5409 = _ctrlsignals_T_273 ? 1'h0 : _ctrlsignals_T_5408; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5410 = _ctrlsignals_T_271 ? 1'h0 : _ctrlsignals_T_5409; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5411 = _ctrlsignals_T_269 ? 1'h0 : _ctrlsignals_T_5410; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5412 = _ctrlsignals_T_267 ? 1'h0 : _ctrlsignals_T_5411; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5413 = _ctrlsignals_T_265 ? 1'h0 : _ctrlsignals_T_5412; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5414 = _ctrlsignals_T_263 ? 1'h0 : _ctrlsignals_T_5413; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5415 = _ctrlsignals_T_261 ? 1'h0 : _ctrlsignals_T_5414; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5416 = _ctrlsignals_T_259 ? 1'h0 : _ctrlsignals_T_5415; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5417 = _ctrlsignals_T_257 ? 1'h0 : _ctrlsignals_T_5416; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5418 = _ctrlsignals_T_255 ? 1'h0 : _ctrlsignals_T_5417; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5419 = _ctrlsignals_T_253 ? 1'h0 : _ctrlsignals_T_5418; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5420 = _ctrlsignals_T_251 ? 1'h0 : _ctrlsignals_T_5419; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5421 = _ctrlsignals_T_249 ? 1'h0 : _ctrlsignals_T_5420; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5422 = _ctrlsignals_T_247 ? 1'h0 : _ctrlsignals_T_5421; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5423 = _ctrlsignals_T_245 ? 1'h0 : _ctrlsignals_T_5422; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5424 = _ctrlsignals_T_243 ? 1'h0 : _ctrlsignals_T_5423; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5425 = _ctrlsignals_T_241 ? 1'h0 : _ctrlsignals_T_5424; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5426 = _ctrlsignals_T_239 ? 1'h0 : _ctrlsignals_T_5425; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5427 = _ctrlsignals_T_237 ? 1'h0 : _ctrlsignals_T_5426; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5428 = _ctrlsignals_T_235 ? 1'h0 : _ctrlsignals_T_5427; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5429 = _ctrlsignals_T_233 ? 1'h0 : _ctrlsignals_T_5428; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5430 = _ctrlsignals_T_231 ? 1'h0 : _ctrlsignals_T_5429; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5431 = _ctrlsignals_T_229 ? 1'h0 : _ctrlsignals_T_5430; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5432 = _ctrlsignals_T_227 ? 1'h0 : _ctrlsignals_T_5431; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5433 = _ctrlsignals_T_225 ? 1'h0 : _ctrlsignals_T_5432; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5434 = _ctrlsignals_T_223 ? 1'h0 : _ctrlsignals_T_5433; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5435 = _ctrlsignals_T_221 ? 1'h0 : _ctrlsignals_T_5434; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5436 = _ctrlsignals_T_219 ? 1'h0 : _ctrlsignals_T_5435; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5437 = _ctrlsignals_T_217 ? 1'h0 : _ctrlsignals_T_5436; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5438 = _ctrlsignals_T_215 ? 1'h0 : _ctrlsignals_T_5437; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5439 = _ctrlsignals_T_213 ? 1'h0 : _ctrlsignals_T_5438; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5440 = _ctrlsignals_T_211 ? 1'h0 : _ctrlsignals_T_5439; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5441 = _ctrlsignals_T_209 ? 1'h0 : _ctrlsignals_T_5440; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5442 = _ctrlsignals_T_207 ? 1'h0 : _ctrlsignals_T_5441; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5443 = _ctrlsignals_T_205 ? 1'h0 : _ctrlsignals_T_5442; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5444 = _ctrlsignals_T_203 ? 1'h0 : _ctrlsignals_T_5443; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5445 = _ctrlsignals_T_201 ? 1'h0 : _ctrlsignals_T_5444; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5446 = _ctrlsignals_T_199 ? 1'h0 : _ctrlsignals_T_5445; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5447 = _ctrlsignals_T_197 ? 1'h0 : _ctrlsignals_T_5446; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5448 = _ctrlsignals_T_195 ? 1'h0 : _ctrlsignals_T_5447; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5449 = _ctrlsignals_T_193 ? 1'h0 : _ctrlsignals_T_5448; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5450 = _ctrlsignals_T_191 ? 1'h0 : _ctrlsignals_T_5449; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5451 = _ctrlsignals_T_189 ? 1'h0 : _ctrlsignals_T_5450; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5452 = _ctrlsignals_T_187 ? 1'h0 : _ctrlsignals_T_5451; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5453 = _ctrlsignals_T_185 ? 1'h0 : _ctrlsignals_T_5452; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5454 = _ctrlsignals_T_183 ? 1'h0 : _ctrlsignals_T_5453; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5455 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_5454; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5456 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_5455; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5457 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_5456; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5458 = _ctrlsignals_T_175 ? 1'h0 : _ctrlsignals_T_5457; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5459 = _ctrlsignals_T_173 ? 1'h0 : _ctrlsignals_T_5458; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5460 = _ctrlsignals_T_171 ? 1'h0 : _ctrlsignals_T_5459; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5461 = _ctrlsignals_T_169 ? 1'h0 : _ctrlsignals_T_5460; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5462 = _ctrlsignals_T_167 ? 1'h0 : _ctrlsignals_T_5461; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5463 = _ctrlsignals_T_165 ? 1'h0 : _ctrlsignals_T_5462; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5464 = _ctrlsignals_T_163 ? 1'h0 : _ctrlsignals_T_5463; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5465 = _ctrlsignals_T_161 ? 1'h0 : _ctrlsignals_T_5464; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5466 = _ctrlsignals_T_159 ? 1'h0 : _ctrlsignals_T_5465; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5467 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_5466; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5468 = _ctrlsignals_T_155 ? 1'h0 : _ctrlsignals_T_5467; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5469 = _ctrlsignals_T_153 ? 1'h0 : _ctrlsignals_T_5468; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5470 = _ctrlsignals_T_151 ? 1'h0 : _ctrlsignals_T_5469; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5471 = _ctrlsignals_T_149 ? 1'h0 : _ctrlsignals_T_5470; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5472 = _ctrlsignals_T_147 ? 1'h0 : _ctrlsignals_T_5471; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5473 = _ctrlsignals_T_145 ? 1'h0 : _ctrlsignals_T_5472; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5474 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_5473; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5475 = _ctrlsignals_T_141 ? 1'h0 : _ctrlsignals_T_5474; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5476 = _ctrlsignals_T_139 ? 1'h0 : _ctrlsignals_T_5475; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5477 = _ctrlsignals_T_137 ? 1'h0 : _ctrlsignals_T_5476; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5478 = _ctrlsignals_T_135 ? 1'h0 : _ctrlsignals_T_5477; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5479 = _ctrlsignals_T_133 ? 1'h0 : _ctrlsignals_T_5478; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5480 = _ctrlsignals_T_131 ? 1'h0 : _ctrlsignals_T_5479; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5481 = _ctrlsignals_T_129 ? 1'h0 : _ctrlsignals_T_5480; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5482 = _ctrlsignals_T_127 ? 1'h0 : _ctrlsignals_T_5481; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5483 = _ctrlsignals_T_125 ? 1'h0 : _ctrlsignals_T_5482; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5484 = _ctrlsignals_T_123 ? 1'h0 : _ctrlsignals_T_5483; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5485 = _ctrlsignals_T_121 ? 1'h0 : _ctrlsignals_T_5484; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5486 = _ctrlsignals_T_119 ? 1'h0 : _ctrlsignals_T_5485; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5487 = _ctrlsignals_T_117 ? 1'h0 : _ctrlsignals_T_5486; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5488 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_5487; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5489 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_5488; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5490 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_5489; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5491 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_5490; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5492 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_5491; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5493 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_5492; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5494 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_5493; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5495 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_5494; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5496 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_5495; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5497 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_5496; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5498 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_5497; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5499 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_5498; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5500 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_5499; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5501 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_5500; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5502 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_5501; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5503 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_5502; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5504 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_5503; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5505 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_5504; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5506 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_5505; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5507 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_5506; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5508 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_5507; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5509 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_5508; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5510 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_5509; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5511 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_5510; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5512 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_5511; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5513 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_5512; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5514 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_5513; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5515 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_5514; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5516 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_5515; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5517 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_5516; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5518 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_5517; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5519 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_5518; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5520 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_5519; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5521 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_5520; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5522 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_5521; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5523 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_5522; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5524 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_5523; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5525 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_5524; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5526 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_5525; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5527 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_5526; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5528 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_5527; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5529 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_5528; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5530 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_5529; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5531 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_5530; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5532 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_5531; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5533 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_5532; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5534 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_5533; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5535 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_5534; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5536 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_5535; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5537 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_5536; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5538 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_5537; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5539 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_5538; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5540 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_5539; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5541 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_5540; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5542 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_5541; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5543 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_5542; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5544 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_5543; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5624 = _ctrlsignals_T_325 ? 1'h0 : _ctrlsignals_T_327 | (_ctrlsignals_T_329 | (_ctrlsignals_T_331
     | (_ctrlsignals_T_333 | (_ctrlsignals_T_335 | (_ctrlsignals_T_337 | (_ctrlsignals_T_339 | (_ctrlsignals_T_341 | (
    _ctrlsignals_T_343 | (_ctrlsignals_T_345 | (_ctrlsignals_T_347 | (_ctrlsignals_T_349 | (_ctrlsignals_T_351 | (
    _ctrlsignals_T_353 | (_ctrlsignals_T_355 | (_ctrlsignals_T_357 | (_ctrlsignals_T_359 | _ctrlsignals_T_361)))))))))))
    ))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5625 = _ctrlsignals_T_323 ? 1'h0 : _ctrlsignals_T_5624; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5626 = _ctrlsignals_T_321 ? 1'h0 : _ctrlsignals_T_5625; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5627 = _ctrlsignals_T_319 ? 1'h0 : _ctrlsignals_T_5626; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5628 = _ctrlsignals_T_317 ? 1'h0 : _ctrlsignals_T_5627; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5629 = _ctrlsignals_T_315 ? 1'h0 : _ctrlsignals_T_5628; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5630 = _ctrlsignals_T_313 ? 1'h0 : _ctrlsignals_T_5629; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5631 = _ctrlsignals_T_311 ? 1'h0 : _ctrlsignals_T_5630; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5632 = _ctrlsignals_T_309 ? 1'h0 : _ctrlsignals_T_5631; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5633 = _ctrlsignals_T_307 ? 1'h0 : _ctrlsignals_T_5632; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5634 = _ctrlsignals_T_305 ? 1'h0 : _ctrlsignals_T_5633; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5635 = _ctrlsignals_T_303 ? 1'h0 : _ctrlsignals_T_5634; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5636 = _ctrlsignals_T_301 ? 1'h0 : _ctrlsignals_T_5635; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5637 = _ctrlsignals_T_299 ? 1'h0 : _ctrlsignals_T_5636; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5638 = _ctrlsignals_T_297 ? 1'h0 : _ctrlsignals_T_5637; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5639 = _ctrlsignals_T_295 ? 1'h0 : _ctrlsignals_T_5638; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5640 = _ctrlsignals_T_293 ? 1'h0 : _ctrlsignals_T_5639; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5641 = _ctrlsignals_T_291 ? 1'h0 : _ctrlsignals_T_5640; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5642 = _ctrlsignals_T_289 ? 1'h0 : _ctrlsignals_T_5641; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5643 = _ctrlsignals_T_287 ? 1'h0 : _ctrlsignals_T_5642; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5644 = _ctrlsignals_T_285 ? 1'h0 : _ctrlsignals_T_5643; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5645 = _ctrlsignals_T_283 ? 1'h0 : _ctrlsignals_T_5644; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5646 = _ctrlsignals_T_281 ? 1'h0 : _ctrlsignals_T_5645; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5647 = _ctrlsignals_T_279 ? 1'h0 : _ctrlsignals_T_5646; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5648 = _ctrlsignals_T_277 ? 1'h0 : _ctrlsignals_T_5647; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5649 = _ctrlsignals_T_275 ? 1'h0 : _ctrlsignals_T_5648; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5650 = _ctrlsignals_T_273 ? 1'h0 : _ctrlsignals_T_5649; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5651 = _ctrlsignals_T_271 ? 1'h0 : _ctrlsignals_T_5650; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5652 = _ctrlsignals_T_269 ? 1'h0 : _ctrlsignals_T_5651; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5653 = _ctrlsignals_T_267 ? 1'h0 : _ctrlsignals_T_5652; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5654 = _ctrlsignals_T_265 ? 1'h0 : _ctrlsignals_T_5653; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5655 = _ctrlsignals_T_263 ? 1'h0 : _ctrlsignals_T_5654; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5656 = _ctrlsignals_T_261 ? 1'h0 : _ctrlsignals_T_5655; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5657 = _ctrlsignals_T_259 ? 1'h0 : _ctrlsignals_T_5656; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5658 = _ctrlsignals_T_257 ? 1'h0 : _ctrlsignals_T_5657; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5659 = _ctrlsignals_T_255 ? 1'h0 : _ctrlsignals_T_5658; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5660 = _ctrlsignals_T_253 ? 1'h0 : _ctrlsignals_T_5659; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5661 = _ctrlsignals_T_251 ? 1'h0 : _ctrlsignals_T_5660; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5662 = _ctrlsignals_T_249 ? 1'h0 : _ctrlsignals_T_5661; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5663 = _ctrlsignals_T_247 ? 1'h0 : _ctrlsignals_T_5662; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5664 = _ctrlsignals_T_245 ? 1'h0 : _ctrlsignals_T_5663; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5665 = _ctrlsignals_T_243 ? 1'h0 : _ctrlsignals_T_5664; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5666 = _ctrlsignals_T_241 ? 1'h0 : _ctrlsignals_T_5665; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5667 = _ctrlsignals_T_239 ? 1'h0 : _ctrlsignals_T_5666; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5668 = _ctrlsignals_T_237 ? 1'h0 : _ctrlsignals_T_5667; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5669 = _ctrlsignals_T_235 ? 1'h0 : _ctrlsignals_T_5668; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5670 = _ctrlsignals_T_233 ? 1'h0 : _ctrlsignals_T_5669; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5671 = _ctrlsignals_T_231 ? 1'h0 : _ctrlsignals_T_5670; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5672 = _ctrlsignals_T_229 ? 1'h0 : _ctrlsignals_T_5671; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5673 = _ctrlsignals_T_227 ? 1'h0 : _ctrlsignals_T_5672; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5674 = _ctrlsignals_T_225 ? 1'h0 : _ctrlsignals_T_5673; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5675 = _ctrlsignals_T_223 ? 1'h0 : _ctrlsignals_T_5674; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5676 = _ctrlsignals_T_221 ? 1'h0 : _ctrlsignals_T_5675; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5677 = _ctrlsignals_T_219 ? 1'h0 : _ctrlsignals_T_5676; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5678 = _ctrlsignals_T_217 ? 1'h0 : _ctrlsignals_T_5677; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5679 = _ctrlsignals_T_215 ? 1'h0 : _ctrlsignals_T_5678; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5680 = _ctrlsignals_T_213 ? 1'h0 : _ctrlsignals_T_5679; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5681 = _ctrlsignals_T_211 ? 1'h0 : _ctrlsignals_T_5680; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5682 = _ctrlsignals_T_209 ? 1'h0 : _ctrlsignals_T_5681; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5683 = _ctrlsignals_T_207 ? 1'h0 : _ctrlsignals_T_5682; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5684 = _ctrlsignals_T_205 ? 1'h0 : _ctrlsignals_T_5683; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5685 = _ctrlsignals_T_203 ? 1'h0 : _ctrlsignals_T_5684; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5686 = _ctrlsignals_T_201 ? 1'h0 : _ctrlsignals_T_5685; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5687 = _ctrlsignals_T_199 ? 1'h0 : _ctrlsignals_T_5686; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5688 = _ctrlsignals_T_197 ? 1'h0 : _ctrlsignals_T_5687; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5689 = _ctrlsignals_T_195 ? 1'h0 : _ctrlsignals_T_5688; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5690 = _ctrlsignals_T_193 ? 1'h0 : _ctrlsignals_T_5689; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5691 = _ctrlsignals_T_191 ? 1'h0 : _ctrlsignals_T_5690; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5692 = _ctrlsignals_T_189 ? 1'h0 : _ctrlsignals_T_5691; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5693 = _ctrlsignals_T_187 ? 1'h0 : _ctrlsignals_T_5692; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5694 = _ctrlsignals_T_185 ? 1'h0 : _ctrlsignals_T_5693; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5695 = _ctrlsignals_T_183 ? 1'h0 : _ctrlsignals_T_5694; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5696 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_5695; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5697 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_5696; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5698 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_5697; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5699 = _ctrlsignals_T_175 ? 1'h0 : _ctrlsignals_T_5698; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5700 = _ctrlsignals_T_173 ? 1'h0 : _ctrlsignals_T_5699; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5701 = _ctrlsignals_T_171 ? 1'h0 : _ctrlsignals_T_5700; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5702 = _ctrlsignals_T_169 ? 1'h0 : _ctrlsignals_T_5701; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5703 = _ctrlsignals_T_167 ? 1'h0 : _ctrlsignals_T_5702; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5704 = _ctrlsignals_T_165 ? 1'h0 : _ctrlsignals_T_5703; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5705 = _ctrlsignals_T_163 ? 1'h0 : _ctrlsignals_T_5704; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5706 = _ctrlsignals_T_161 ? 1'h0 : _ctrlsignals_T_5705; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5707 = _ctrlsignals_T_159 ? 1'h0 : _ctrlsignals_T_5706; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5708 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_5707; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5709 = _ctrlsignals_T_155 ? 1'h0 : _ctrlsignals_T_5708; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5710 = _ctrlsignals_T_153 ? 1'h0 : _ctrlsignals_T_5709; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5711 = _ctrlsignals_T_151 ? 1'h0 : _ctrlsignals_T_5710; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5712 = _ctrlsignals_T_149 ? 1'h0 : _ctrlsignals_T_5711; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5713 = _ctrlsignals_T_147 ? 1'h0 : _ctrlsignals_T_5712; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5714 = _ctrlsignals_T_145 ? 1'h0 : _ctrlsignals_T_5713; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5715 = _ctrlsignals_T_143 ? 1'h0 : _ctrlsignals_T_5714; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5716 = _ctrlsignals_T_141 ? 1'h0 : _ctrlsignals_T_5715; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5717 = _ctrlsignals_T_139 ? 1'h0 : _ctrlsignals_T_5716; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5718 = _ctrlsignals_T_137 ? 1'h0 : _ctrlsignals_T_5717; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5719 = _ctrlsignals_T_135 ? 1'h0 : _ctrlsignals_T_5718; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5720 = _ctrlsignals_T_133 ? 1'h0 : _ctrlsignals_T_5719; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5721 = _ctrlsignals_T_131 ? 1'h0 : _ctrlsignals_T_5720; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5722 = _ctrlsignals_T_129 ? 1'h0 : _ctrlsignals_T_5721; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5723 = _ctrlsignals_T_127 ? 1'h0 : _ctrlsignals_T_5722; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5724 = _ctrlsignals_T_125 ? 1'h0 : _ctrlsignals_T_5723; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5725 = _ctrlsignals_T_123 ? 1'h0 : _ctrlsignals_T_5724; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5726 = _ctrlsignals_T_121 ? 1'h0 : _ctrlsignals_T_5725; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5727 = _ctrlsignals_T_119 ? 1'h0 : _ctrlsignals_T_5726; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5728 = _ctrlsignals_T_117 ? 1'h0 : _ctrlsignals_T_5727; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5729 = _ctrlsignals_T_115 ? 1'h0 : _ctrlsignals_T_5728; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5730 = _ctrlsignals_T_113 ? 1'h0 : _ctrlsignals_T_5729; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5731 = _ctrlsignals_T_111 ? 1'h0 : _ctrlsignals_T_5730; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5732 = _ctrlsignals_T_109 ? 1'h0 : _ctrlsignals_T_5731; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5733 = _ctrlsignals_T_107 ? 1'h0 : _ctrlsignals_T_5732; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5734 = _ctrlsignals_T_105 ? 1'h0 : _ctrlsignals_T_5733; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5735 = _ctrlsignals_T_103 ? 1'h0 : _ctrlsignals_T_5734; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5736 = _ctrlsignals_T_101 ? 1'h0 : _ctrlsignals_T_5735; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5737 = _ctrlsignals_T_99 ? 1'h0 : _ctrlsignals_T_5736; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5738 = _ctrlsignals_T_97 ? 1'h0 : _ctrlsignals_T_5737; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5739 = _ctrlsignals_T_95 ? 1'h0 : _ctrlsignals_T_5738; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5740 = _ctrlsignals_T_93 ? 1'h0 : _ctrlsignals_T_5739; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5741 = _ctrlsignals_T_91 ? 1'h0 : _ctrlsignals_T_5740; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5742 = _ctrlsignals_T_89 ? 1'h0 : _ctrlsignals_T_5741; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5743 = _ctrlsignals_T_87 ? 1'h0 : _ctrlsignals_T_5742; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5744 = _ctrlsignals_T_85 ? 1'h0 : _ctrlsignals_T_5743; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5745 = _ctrlsignals_T_83 ? 1'h0 : _ctrlsignals_T_5744; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5746 = _ctrlsignals_T_81 ? 1'h0 : _ctrlsignals_T_5745; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5747 = _ctrlsignals_T_79 ? 1'h0 : _ctrlsignals_T_5746; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5748 = _ctrlsignals_T_77 ? 1'h0 : _ctrlsignals_T_5747; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5749 = _ctrlsignals_T_75 ? 1'h0 : _ctrlsignals_T_5748; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5750 = _ctrlsignals_T_73 ? 1'h0 : _ctrlsignals_T_5749; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5751 = _ctrlsignals_T_71 ? 1'h0 : _ctrlsignals_T_5750; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5752 = _ctrlsignals_T_69 ? 1'h0 : _ctrlsignals_T_5751; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5753 = _ctrlsignals_T_67 ? 1'h0 : _ctrlsignals_T_5752; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5754 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_5753; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5755 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_5754; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5756 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_5755; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5757 = _ctrlsignals_T_59 ? 1'h0 : _ctrlsignals_T_5756; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5758 = _ctrlsignals_T_57 ? 1'h0 : _ctrlsignals_T_5757; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5759 = _ctrlsignals_T_55 ? 1'h0 : _ctrlsignals_T_5758; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5760 = _ctrlsignals_T_53 ? 1'h0 : _ctrlsignals_T_5759; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5761 = _ctrlsignals_T_51 ? 1'h0 : _ctrlsignals_T_5760; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5762 = _ctrlsignals_T_49 ? 1'h0 : _ctrlsignals_T_5761; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5763 = _ctrlsignals_T_47 ? 1'h0 : _ctrlsignals_T_5762; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5764 = _ctrlsignals_T_45 ? 1'h0 : _ctrlsignals_T_5763; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5765 = _ctrlsignals_T_43 ? 1'h0 : _ctrlsignals_T_5764; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5766 = _ctrlsignals_T_41 ? 1'h0 : _ctrlsignals_T_5765; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5767 = _ctrlsignals_T_39 ? 1'h0 : _ctrlsignals_T_5766; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5768 = _ctrlsignals_T_37 ? 1'h0 : _ctrlsignals_T_5767; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5769 = _ctrlsignals_T_35 ? 1'h0 : _ctrlsignals_T_5768; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5770 = _ctrlsignals_T_33 ? 1'h0 : _ctrlsignals_T_5769; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5771 = _ctrlsignals_T_31 ? 1'h0 : _ctrlsignals_T_5770; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5772 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_5771; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5773 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_5772; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5774 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_5773; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5775 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_5774; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5776 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_5775; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5777 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_5776; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5778 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_5777; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5779 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_5778; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5780 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_5779; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5781 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_5780; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5782 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_5781; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5783 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_5782; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5784 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_5783; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5785 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_5784; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5790 = _ctrlsignals_T_475 ? 1'h0 : _ctrlsignals_T_477; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5791 = _ctrlsignals_T_473 ? 1'h0 : _ctrlsignals_T_5790; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5792 = _ctrlsignals_T_471 ? 1'h0 : _ctrlsignals_T_5791; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5793 = _ctrlsignals_T_469 ? 1'h0 : _ctrlsignals_T_5792; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5794 = _ctrlsignals_T_467 ? 1'h0 : _ctrlsignals_T_5793; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5795 = _ctrlsignals_T_465 ? 1'h0 : _ctrlsignals_T_5794; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5796 = _ctrlsignals_T_463 ? 1'h0 : _ctrlsignals_T_5795; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5797 = _ctrlsignals_T_461 ? 1'h0 : _ctrlsignals_T_5796; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5798 = _ctrlsignals_T_459 ? 1'h0 : _ctrlsignals_T_5797; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5799 = _ctrlsignals_T_445 ? 1'h0 : _ctrlsignals_T_5798; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5800 = _ctrlsignals_T_443 ? 1'h0 : _ctrlsignals_T_5799; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5801 = _ctrlsignals_T_453 ? 1'h0 : _ctrlsignals_T_5800; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5802 = _ctrlsignals_T_451 ? 1'h0 : _ctrlsignals_T_5801; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5803 = _ctrlsignals_T_449 ? 1'h0 : _ctrlsignals_T_5802; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5804 = _ctrlsignals_T_447 ? 1'h0 : _ctrlsignals_T_5803; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5805 = _ctrlsignals_T_445 ? 1'h0 : _ctrlsignals_T_5804; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5806 = _ctrlsignals_T_443 ? 1'h0 : _ctrlsignals_T_5805; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5807 = _ctrlsignals_T_441 ? 1'h0 : _ctrlsignals_T_5806; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5808 = _ctrlsignals_T_439 ? 1'h0 : _ctrlsignals_T_5807; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5809 = _ctrlsignals_T_437 ? 1'h0 : _ctrlsignals_T_5808; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5810 = _ctrlsignals_T_435 ? 1'h0 : _ctrlsignals_T_5809; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5811 = _ctrlsignals_T_433 ? 1'h0 : _ctrlsignals_T_5810; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5812 = _ctrlsignals_T_431 ? 1'h0 : _ctrlsignals_T_5811; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5813 = _ctrlsignals_T_429 ? 1'h0 : _ctrlsignals_T_5812; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5814 = _ctrlsignals_T_427 ? 1'h0 : _ctrlsignals_T_5813; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5815 = _ctrlsignals_T_425 ? 1'h0 : _ctrlsignals_T_5814; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5816 = _ctrlsignals_T_423 ? 1'h0 : _ctrlsignals_T_5815; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5817 = _ctrlsignals_T_421 ? 1'h0 : _ctrlsignals_T_5816; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5818 = _ctrlsignals_T_419 ? 1'h0 : _ctrlsignals_T_5817; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5819 = _ctrlsignals_T_417 ? 1'h0 : _ctrlsignals_T_5818; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5820 = _ctrlsignals_T_415 ? 1'h0 : _ctrlsignals_T_5819; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5821 = _ctrlsignals_T_413 ? 1'h0 : _ctrlsignals_T_5820; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5822 = _ctrlsignals_T_411 ? 1'h0 : _ctrlsignals_T_5821; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5823 = _ctrlsignals_T_409 ? 1'h0 : _ctrlsignals_T_5822; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5824 = _ctrlsignals_T_407 ? 1'h0 : _ctrlsignals_T_5823; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5825 = _ctrlsignals_T_405 ? 1'h0 : _ctrlsignals_T_5824; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5826 = _ctrlsignals_T_403 ? 1'h0 : _ctrlsignals_T_5825; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5827 = _ctrlsignals_T_401 ? 1'h0 : _ctrlsignals_T_5826; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5828 = _ctrlsignals_T_399 ? 1'h0 : _ctrlsignals_T_5827; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5829 = _ctrlsignals_T_397 ? 1'h0 : _ctrlsignals_T_5828; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5830 = _ctrlsignals_T_395 ? 1'h0 : _ctrlsignals_T_5829; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5831 = _ctrlsignals_T_393 ? 1'h0 : _ctrlsignals_T_5830; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5832 = _ctrlsignals_T_391 ? 1'h0 : _ctrlsignals_T_5831; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5833 = _ctrlsignals_T_389 ? 1'h0 : _ctrlsignals_T_5832; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5834 = _ctrlsignals_T_387 ? 1'h0 : _ctrlsignals_T_5833; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5835 = _ctrlsignals_T_385 ? 1'h0 : _ctrlsignals_T_5834; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5836 = _ctrlsignals_T_383 ? 1'h0 : _ctrlsignals_T_5835; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5837 = _ctrlsignals_T_381 ? 1'h0 : _ctrlsignals_T_5836; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5838 = _ctrlsignals_T_379 ? 1'h0 : _ctrlsignals_T_5837; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5839 = _ctrlsignals_T_377 ? 1'h0 : _ctrlsignals_T_5838; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5840 = _ctrlsignals_T_375 ? 1'h0 : _ctrlsignals_T_5839; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5841 = _ctrlsignals_T_373 ? 1'h0 : _ctrlsignals_T_5840; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5842 = _ctrlsignals_T_371 ? 1'h0 : _ctrlsignals_T_5841; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5843 = _ctrlsignals_T_369 ? 1'h0 : _ctrlsignals_T_5842; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5844 = _ctrlsignals_T_367 ? 1'h0 : _ctrlsignals_T_5843; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5845 = _ctrlsignals_T_365 ? 1'h0 : _ctrlsignals_T_5844; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5846 = _ctrlsignals_T_363 ? 1'h0 : _ctrlsignals_T_5845; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5847 = _ctrlsignals_T_361 ? 1'h0 : _ctrlsignals_T_5846; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5848 = _ctrlsignals_T_359 ? 1'h0 : _ctrlsignals_T_5847; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5849 = _ctrlsignals_T_357 ? 1'h0 : _ctrlsignals_T_5848; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5850 = _ctrlsignals_T_355 ? 1'h0 : _ctrlsignals_T_5849; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5851 = _ctrlsignals_T_353 ? 1'h0 : _ctrlsignals_T_5850; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5852 = _ctrlsignals_T_351 ? 1'h0 : _ctrlsignals_T_5851; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5853 = _ctrlsignals_T_349 ? 1'h0 : _ctrlsignals_T_5852; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5854 = _ctrlsignals_T_347 ? 1'h0 : _ctrlsignals_T_5853; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5855 = _ctrlsignals_T_345 ? 1'h0 : _ctrlsignals_T_5854; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5856 = _ctrlsignals_T_343 ? 1'h0 : _ctrlsignals_T_5855; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5857 = _ctrlsignals_T_341 ? 1'h0 : _ctrlsignals_T_5856; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5858 = _ctrlsignals_T_339 ? 1'h0 : _ctrlsignals_T_5857; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5859 = _ctrlsignals_T_337 ? 1'h0 : _ctrlsignals_T_5858; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5860 = _ctrlsignals_T_335 ? 1'h0 : _ctrlsignals_T_5859; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5861 = _ctrlsignals_T_333 ? 1'h0 : _ctrlsignals_T_5860; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5862 = _ctrlsignals_T_331 ? 1'h0 : _ctrlsignals_T_5861; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5863 = _ctrlsignals_T_329 ? 1'h0 : _ctrlsignals_T_5862; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5864 = _ctrlsignals_T_327 ? 1'h0 : _ctrlsignals_T_5863; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5865 = _ctrlsignals_T_325 ? 1'h0 : _ctrlsignals_T_5864; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5866 = _ctrlsignals_T_323 ? 1'h0 : _ctrlsignals_T_5865; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5867 = _ctrlsignals_T_321 ? 1'h0 : _ctrlsignals_T_5866; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5868 = _ctrlsignals_T_319 ? 1'h0 : _ctrlsignals_T_5867; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5869 = _ctrlsignals_T_317 ? 1'h0 : _ctrlsignals_T_5868; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5870 = _ctrlsignals_T_315 ? 1'h0 : _ctrlsignals_T_5869; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5871 = _ctrlsignals_T_313 ? 1'h0 : _ctrlsignals_T_5870; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5872 = _ctrlsignals_T_311 ? 1'h0 : _ctrlsignals_T_5871; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5873 = _ctrlsignals_T_309 ? 1'h0 : _ctrlsignals_T_5872; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5874 = _ctrlsignals_T_307 ? 1'h0 : _ctrlsignals_T_5873; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5875 = _ctrlsignals_T_305 ? 1'h0 : _ctrlsignals_T_5874; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5876 = _ctrlsignals_T_303 ? 1'h0 : _ctrlsignals_T_5875; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5877 = _ctrlsignals_T_301 ? 1'h0 : _ctrlsignals_T_5876; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5878 = _ctrlsignals_T_299 ? 1'h0 : _ctrlsignals_T_5877; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5879 = _ctrlsignals_T_297 ? 1'h0 : _ctrlsignals_T_5878; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5880 = _ctrlsignals_T_295 ? 1'h0 : _ctrlsignals_T_5879; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5881 = _ctrlsignals_T_293 ? 1'h0 : _ctrlsignals_T_5880; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5882 = _ctrlsignals_T_291 ? 1'h0 : _ctrlsignals_T_5881; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5883 = _ctrlsignals_T_289 ? 1'h0 : _ctrlsignals_T_5882; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5884 = _ctrlsignals_T_287 ? 1'h0 : _ctrlsignals_T_5883; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5885 = _ctrlsignals_T_285 ? 1'h0 : _ctrlsignals_T_5884; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5886 = _ctrlsignals_T_283 ? 1'h0 : _ctrlsignals_T_5885; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5887 = _ctrlsignals_T_281 ? 1'h0 : _ctrlsignals_T_5886; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5888 = _ctrlsignals_T_279 ? 1'h0 : _ctrlsignals_T_5887; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5889 = _ctrlsignals_T_277 ? 1'h0 : _ctrlsignals_T_5888; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5890 = _ctrlsignals_T_275 ? 1'h0 : _ctrlsignals_T_5889; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5891 = _ctrlsignals_T_273 ? 1'h0 : _ctrlsignals_T_5890; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5892 = _ctrlsignals_T_271 ? 1'h0 : _ctrlsignals_T_5891; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5893 = _ctrlsignals_T_269 ? 1'h0 : _ctrlsignals_T_5892; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5894 = _ctrlsignals_T_267 ? 1'h0 : _ctrlsignals_T_5893; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5895 = _ctrlsignals_T_265 ? 1'h0 : _ctrlsignals_T_5894; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5896 = _ctrlsignals_T_263 ? 1'h0 : _ctrlsignals_T_5895; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5897 = _ctrlsignals_T_261 ? 1'h0 : _ctrlsignals_T_5896; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5898 = _ctrlsignals_T_259 ? 1'h0 : _ctrlsignals_T_5897; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5899 = _ctrlsignals_T_257 ? 1'h0 : _ctrlsignals_T_5898; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5900 = _ctrlsignals_T_255 ? 1'h0 : _ctrlsignals_T_5899; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5901 = _ctrlsignals_T_253 ? 1'h0 : _ctrlsignals_T_5900; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5902 = _ctrlsignals_T_251 ? 1'h0 : _ctrlsignals_T_5901; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5903 = _ctrlsignals_T_249 ? 1'h0 : _ctrlsignals_T_5902; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5904 = _ctrlsignals_T_247 ? 1'h0 : _ctrlsignals_T_5903; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5905 = _ctrlsignals_T_245 ? 1'h0 : _ctrlsignals_T_5904; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5906 = _ctrlsignals_T_243 ? 1'h0 : _ctrlsignals_T_5905; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5907 = _ctrlsignals_T_241 ? 1'h0 : _ctrlsignals_T_5906; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5908 = _ctrlsignals_T_239 ? 1'h0 : _ctrlsignals_T_5907; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5909 = _ctrlsignals_T_237 ? 1'h0 : _ctrlsignals_T_5908; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5910 = _ctrlsignals_T_235 ? 1'h0 : _ctrlsignals_T_5909; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5911 = _ctrlsignals_T_233 ? 1'h0 : _ctrlsignals_T_5910; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5912 = _ctrlsignals_T_231 ? 1'h0 : _ctrlsignals_T_5911; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5913 = _ctrlsignals_T_229 ? 1'h0 : _ctrlsignals_T_5912; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5914 = _ctrlsignals_T_227 ? 1'h0 : _ctrlsignals_T_5913; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5915 = _ctrlsignals_T_225 ? 1'h0 : _ctrlsignals_T_5914; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5916 = _ctrlsignals_T_223 ? 1'h0 : _ctrlsignals_T_5915; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5917 = _ctrlsignals_T_221 ? 1'h0 : _ctrlsignals_T_5916; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5918 = _ctrlsignals_T_219 ? 1'h0 : _ctrlsignals_T_5917; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5919 = _ctrlsignals_T_217 ? 1'h0 : _ctrlsignals_T_5918; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5920 = _ctrlsignals_T_215 ? 1'h0 : _ctrlsignals_T_5919; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5921 = _ctrlsignals_T_213 ? 1'h0 : _ctrlsignals_T_5920; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5922 = _ctrlsignals_T_211 ? 1'h0 : _ctrlsignals_T_5921; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5923 = _ctrlsignals_T_209 ? 1'h0 : _ctrlsignals_T_5922; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5924 = _ctrlsignals_T_207 ? 1'h0 : _ctrlsignals_T_5923; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5925 = _ctrlsignals_T_205 ? 1'h0 : _ctrlsignals_T_5924; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5926 = _ctrlsignals_T_203 ? 1'h0 : _ctrlsignals_T_5925; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5927 = _ctrlsignals_T_201 ? 1'h0 : _ctrlsignals_T_5926; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5928 = _ctrlsignals_T_199 ? 1'h0 : _ctrlsignals_T_5927; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5929 = _ctrlsignals_T_197 ? 1'h0 : _ctrlsignals_T_5928; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5930 = _ctrlsignals_T_195 ? 1'h0 : _ctrlsignals_T_5929; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5931 = _ctrlsignals_T_193 ? 1'h0 : _ctrlsignals_T_5930; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5932 = _ctrlsignals_T_191 ? 1'h0 : _ctrlsignals_T_5931; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5933 = _ctrlsignals_T_189 ? 1'h0 : _ctrlsignals_T_5932; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5934 = _ctrlsignals_T_187 ? 1'h0 : _ctrlsignals_T_5933; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5935 = _ctrlsignals_T_185 ? 1'h0 : _ctrlsignals_T_5934; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5936 = _ctrlsignals_T_183 ? 1'h0 : _ctrlsignals_T_5935; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5937 = _ctrlsignals_T_181 ? 1'h0 : _ctrlsignals_T_5936; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5938 = _ctrlsignals_T_179 ? 1'h0 : _ctrlsignals_T_5937; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5939 = _ctrlsignals_T_177 ? 1'h0 : _ctrlsignals_T_5938; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5940 = _ctrlsignals_T_175 ? 1'h0 : _ctrlsignals_T_5939; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5941 = _ctrlsignals_T_173 ? 1'h0 : _ctrlsignals_T_5940; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5942 = _ctrlsignals_T_171 ? 1'h0 : _ctrlsignals_T_5941; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5972 = _ctrlsignals_T_111 | (_ctrlsignals_T_113 | (_ctrlsignals_T_115 | (_ctrlsignals_T_117 | (
    _ctrlsignals_T_119 | (_ctrlsignals_T_121 | (_ctrlsignals_T_123 | (_ctrlsignals_T_125 | (_ctrlsignals_T_127 | (
    _ctrlsignals_T_129 | (_ctrlsignals_T_131 | (_ctrlsignals_T_133 | (_ctrlsignals_T_135 | (_ctrlsignals_T_137 | (
    _ctrlsignals_T_139 | (_ctrlsignals_T_141 | (_ctrlsignals_T_143 | (_ctrlsignals_T_145 | (_ctrlsignals_T_147 | (
    _ctrlsignals_T_149 | (_ctrlsignals_T_151 | (_ctrlsignals_T_153 | (_ctrlsignals_T_155 | (_ctrlsignals_T_143 | (
    _ctrlsignals_T_159 | (_ctrlsignals_T_161 | (_ctrlsignals_T_163 | (_ctrlsignals_T_165 | (_ctrlsignals_T_167 | (
    _ctrlsignals_T_169 | _ctrlsignals_T_5942))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5995 = _ctrlsignals_T_65 ? 1'h0 : _ctrlsignals_T_67 | (_ctrlsignals_T_69 | (_ctrlsignals_T_71 | (
    _ctrlsignals_T_73 | (_ctrlsignals_T_75 | (_ctrlsignals_T_77 | (_ctrlsignals_T_79 | (_ctrlsignals_T_81 | (
    _ctrlsignals_T_83 | (_ctrlsignals_T_85 | (_ctrlsignals_T_87 | (_ctrlsignals_T_89 | (_ctrlsignals_T_91 | (
    _ctrlsignals_T_93 | (_ctrlsignals_T_95 | (_ctrlsignals_T_97 | (_ctrlsignals_T_99 | (_ctrlsignals_T_101 | (
    _ctrlsignals_T_103 | (_ctrlsignals_T_105 | (_ctrlsignals_T_107 | (_ctrlsignals_T_109 | _ctrlsignals_T_5972))))))))))
    ))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5996 = _ctrlsignals_T_63 ? 1'h0 : _ctrlsignals_T_5995; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_5997 = _ctrlsignals_T_61 ? 1'h0 : _ctrlsignals_T_5996; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6013 = _ctrlsignals_T_29 ? 1'h0 : _ctrlsignals_T_31 | (_ctrlsignals_T_33 | (_ctrlsignals_T_35 | (
    _ctrlsignals_T_37 | (_ctrlsignals_T_39 | (_ctrlsignals_T_41 | (_ctrlsignals_T_43 | (_ctrlsignals_T_45 | (
    _ctrlsignals_T_47 | (_ctrlsignals_T_49 | (_ctrlsignals_T_51 | (_ctrlsignals_T_53 | (_ctrlsignals_T_55 | (
    _ctrlsignals_T_57 | (_ctrlsignals_T_59 | _ctrlsignals_T_5997)))))))))))))); // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6014 = _ctrlsignals_T_27 ? 1'h0 : _ctrlsignals_T_6013; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6015 = _ctrlsignals_T_25 ? 1'h0 : _ctrlsignals_T_6014; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6016 = _ctrlsignals_T_23 ? 1'h0 : _ctrlsignals_T_6015; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6017 = _ctrlsignals_T_21 ? 1'h0 : _ctrlsignals_T_6016; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6018 = _ctrlsignals_T_19 ? 1'h0 : _ctrlsignals_T_6017; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6019 = _ctrlsignals_T_17 ? 1'h0 : _ctrlsignals_T_6018; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6020 = _ctrlsignals_T_15 ? 1'h0 : _ctrlsignals_T_6019; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6021 = _ctrlsignals_T_13 ? 1'h0 : _ctrlsignals_T_6020; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6022 = _ctrlsignals_T_11 ? 1'h0 : _ctrlsignals_T_6021; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6023 = _ctrlsignals_T_9 ? 1'h0 : _ctrlsignals_T_6022; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6024 = _ctrlsignals_T_7 ? 1'h0 : _ctrlsignals_T_6023; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6025 = _ctrlsignals_T_5 ? 1'h0 : _ctrlsignals_T_6024; // @[Lookup.scala 34:39]
  wire  _ctrlsignals_T_6026 = _ctrlsignals_T_3 ? 1'h0 : _ctrlsignals_T_6025; // @[Lookup.scala 34:39]
  assign io_control_inst = io_inst; // @[DecodeUnit.scala 411:18]
  assign io_control_wid = io_wid; // @[DecodeUnit.scala 412:17]
  assign io_control_fp = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_965; // @[Lookup.scala 34:39]
  assign io_control_branch = _ctrlsignals_T_1 ? 2'h1 : _ctrlsignals_T_1447; // @[Lookup.scala 34:39]
  assign io_control_simt_stack = _ctrlsignals_T_1 | (_ctrlsignals_T_3 | (_ctrlsignals_T_5 | (_ctrlsignals_T_7 | (
    _ctrlsignals_T_9 | (_ctrlsignals_T_11 | _ctrlsignals_T_13))))); // @[Lookup.scala 34:39]
  assign io_control_simt_stack_op = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_1929; // @[Lookup.scala 34:39]
  assign io_control_barrier = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_1206; // @[Lookup.scala 34:39]
  assign io_control_csr = _ctrlsignals_T_1 ? 2'h0 : _ctrlsignals_T_2170; // @[Lookup.scala 34:39]
  assign io_control_reverse = _ctrlsignals_T_1 | (_ctrlsignals_T_3 | (_ctrlsignals_T_5 | (_ctrlsignals_T_7 | (
    _ctrlsignals_T_9 | (_ctrlsignals_T_11 | _ctrlsignals_T_2406))))); // @[Lookup.scala 34:39]
  assign io_control_sel_alu2 = _ctrlsignals_T_1 ? 2'h2 : _ctrlsignals_T_2893; // @[Lookup.scala 34:39]
  assign io_control_sel_alu1 = _ctrlsignals_T_1 ? 2'h2 : _ctrlsignals_T_3134; // @[Lookup.scala 34:39]
  assign io_control_isvec = _ctrlsignals_T_1 | (_ctrlsignals_T_3 | (_ctrlsignals_T_5 | (_ctrlsignals_T_7 | (
    _ctrlsignals_T_9 | (_ctrlsignals_T_11 | (_ctrlsignals_T_13 | _ctrlsignals_T_718)))))); // @[Lookup.scala 34:39]
  assign io_control_sel_alu3 = _ctrlsignals_T_1 ? 2'h0 : _ctrlsignals_T_2652; // @[Lookup.scala 34:39]
  assign io_control_mask = (~io_inst[25] | io_control_alu_fn == 6'h13) & io_control_isvec & ~(|io_control_branch); // @[DecodeUnit.scala 424:115]
  assign io_control_sel_imm = _ctrlsignals_T_1 ? 3'h2 : _ctrlsignals_T_3375; // @[Lookup.scala 34:39]
  assign io_control_mem_unsigned = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_4580; // @[Lookup.scala 34:39]
  assign io_control_alu_fn = _ctrlsignals_T_1 ? 6'h3 : _ctrlsignals_T_3857; // @[Lookup.scala 34:39]
  assign io_control_mem = |io_control_mem_cmd; // @[DecodeUnit.scala 430:38]
  assign io_control_mem_cmd = _ctrlsignals_T_1 ? 2'h0 : _ctrlsignals_T_4339; // @[Lookup.scala 34:39]
  assign io_control_mop = io_inst[27:26]; // @[DecodeUnit.scala 414:26]
  assign io_control_reg_idx1 = io_inst[19:15]; // @[DecodeUnit.scala 439:31]
  assign io_control_reg_idx2 = io_inst[24:20]; // @[DecodeUnit.scala 440:31]
  assign io_control_reg_idx3 = io_control_fp & ~io_control_isvec ? io_inst[31:27] : io_inst[11:7]; // @[DecodeUnit.scala 441:27]
  assign io_control_reg_idxw = io_inst[11:7]; // @[DecodeUnit.scala 442:31]
  assign io_control_wfd = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_5303; // @[Lookup.scala 34:39]
  assign io_control_fence = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_4821; // @[Lookup.scala 34:39]
  assign io_control_sfu = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_5062; // @[Lookup.scala 34:39]
  assign io_control_readmask = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_5544; // @[Lookup.scala 34:39]
  assign io_control_writemask = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_5785; // @[Lookup.scala 34:39]
  assign io_control_wxd = _ctrlsignals_T_1 ? 1'h0 : _ctrlsignals_T_6026; // @[Lookup.scala 34:39]
  assign io_control_pc = io_pc; // @[DecodeUnit.scala 413:16]
endmodule
module FloatRegFile(
  input         clock,
  output [31:0] io_v0_0,
  output [31:0] io_rs1_0,
  output [31:0] io_rs1_1,
  output [31:0] io_rs1_2,
  output [31:0] io_rs1_3,
  output [31:0] io_rs1_4,
  output [31:0] io_rs1_5,
  output [31:0] io_rs1_6,
  output [31:0] io_rs1_7,
  output [31:0] io_rs2_0,
  output [31:0] io_rs2_1,
  output [31:0] io_rs2_2,
  output [31:0] io_rs2_3,
  output [31:0] io_rs2_4,
  output [31:0] io_rs2_5,
  output [31:0] io_rs2_6,
  output [31:0] io_rs2_7,
  output [31:0] io_rs3_0,
  output [31:0] io_rs3_1,
  output [31:0] io_rs3_2,
  output [31:0] io_rs3_3,
  output [31:0] io_rs3_4,
  output [31:0] io_rs3_5,
  output [31:0] io_rs3_6,
  output [31:0] io_rs3_7,
  input  [4:0]  io_rs1idx,
  input  [4:0]  io_rs2idx,
  input  [4:0]  io_rs3idx,
  input  [31:0] io_rd_0,
  input  [31:0] io_rd_1,
  input  [31:0] io_rd_2,
  input  [31:0] io_rd_3,
  input  [31:0] io_rd_4,
  input  [31:0] io_rd_5,
  input  [31:0] io_rd_6,
  input  [31:0] io_rd_7,
  input  [4:0]  io_rdidx,
  input         io_rdwen,
  input         io_rdwmask_0,
  input         io_rdwmask_1,
  input         io_rdwmask_2,
  input         io_rdwmask_3,
  input         io_rdwmask_4,
  input         io_rdwmask_5,
  input         io_rdwmask_6,
  input         io_rdwmask_7
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] regs_0 [0:31]; // @[regfile.scala 49:17]
  wire  regs_0_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_0_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_0_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_0_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_0_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_0_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_0_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_0_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_0_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_0_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_0_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_0_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_0_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_0_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_0_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_0_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_1 [0:31]; // @[regfile.scala 49:17]
  wire  regs_1_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_1_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_1_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_1_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_1_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_1_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_1_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_1_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_1_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_1_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_1_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_1_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_1_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_1_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_1_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_1_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_2 [0:31]; // @[regfile.scala 49:17]
  wire  regs_2_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_2_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_2_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_2_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_2_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_2_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_2_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_2_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_2_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_2_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_2_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_2_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_2_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_2_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_2_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_2_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_3 [0:31]; // @[regfile.scala 49:17]
  wire  regs_3_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_3_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_3_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_3_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_3_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_3_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_3_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_3_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_3_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_3_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_3_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_3_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_3_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_3_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_3_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_3_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_4 [0:31]; // @[regfile.scala 49:17]
  wire  regs_4_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_4_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_4_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_4_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_4_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_4_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_4_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_4_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_4_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_4_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_4_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_4_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_4_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_4_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_4_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_4_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_5 [0:31]; // @[regfile.scala 49:17]
  wire  regs_5_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_5_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_5_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_5_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_5_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_5_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_5_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_5_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_5_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_5_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_5_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_5_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_5_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_5_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_5_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_5_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_6 [0:31]; // @[regfile.scala 49:17]
  wire  regs_6_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_6_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_6_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_6_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_6_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_6_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_6_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_6_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_6_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_6_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_6_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_6_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_6_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_6_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_6_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_6_MPORT_4_en; // @[regfile.scala 49:17]
  reg [31:0] regs_7 [0:31]; // @[regfile.scala 49:17]
  wire  regs_7_MPORT_en; // @[regfile.scala 49:17]
  wire [4:0] regs_7_MPORT_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_7_MPORT_data; // @[regfile.scala 49:17]
  wire  regs_7_MPORT_1_en; // @[regfile.scala 49:17]
  wire [4:0] regs_7_MPORT_1_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_7_MPORT_1_data; // @[regfile.scala 49:17]
  wire  regs_7_MPORT_2_en; // @[regfile.scala 49:17]
  wire [4:0] regs_7_MPORT_2_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_7_MPORT_2_data; // @[regfile.scala 49:17]
  wire  regs_7_MPORT_3_en; // @[regfile.scala 49:17]
  wire [4:0] regs_7_MPORT_3_addr; // @[regfile.scala 49:17]
  wire [31:0] regs_7_MPORT_3_data; // @[regfile.scala 49:17]
  wire [31:0] regs_7_MPORT_4_data; // @[regfile.scala 49:17]
  wire [4:0] regs_7_MPORT_4_addr; // @[regfile.scala 49:17]
  wire  regs_7_MPORT_4_mask; // @[regfile.scala 49:17]
  wire  regs_7_MPORT_4_en; // @[regfile.scala 49:17]
  assign regs_0_MPORT_en = 1'h1;
  assign regs_0_MPORT_addr = io_rs1idx;
  assign regs_0_MPORT_data = regs_0[regs_0_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_0_MPORT_1_en = 1'h1;
  assign regs_0_MPORT_1_addr = io_rs2idx;
  assign regs_0_MPORT_1_data = regs_0[regs_0_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_0_MPORT_2_en = 1'h1;
  assign regs_0_MPORT_2_addr = io_rs3idx;
  assign regs_0_MPORT_2_data = regs_0[regs_0_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_0_MPORT_3_en = 1'h1;
  assign regs_0_MPORT_3_addr = 5'h0;
  assign regs_0_MPORT_3_data = regs_0[regs_0_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_0_MPORT_4_data = io_rd_0;
  assign regs_0_MPORT_4_addr = io_rdidx;
  assign regs_0_MPORT_4_mask = io_rdwmask_0;
  assign regs_0_MPORT_4_en = io_rdwen;
  assign regs_1_MPORT_en = 1'h1;
  assign regs_1_MPORT_addr = io_rs1idx;
  assign regs_1_MPORT_data = regs_1[regs_1_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_1_MPORT_1_en = 1'h1;
  assign regs_1_MPORT_1_addr = io_rs2idx;
  assign regs_1_MPORT_1_data = regs_1[regs_1_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_1_MPORT_2_en = 1'h1;
  assign regs_1_MPORT_2_addr = io_rs3idx;
  assign regs_1_MPORT_2_data = regs_1[regs_1_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_1_MPORT_3_en = 1'h1;
  assign regs_1_MPORT_3_addr = 5'h0;
  assign regs_1_MPORT_3_data = regs_1[regs_1_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_1_MPORT_4_data = io_rd_1;
  assign regs_1_MPORT_4_addr = io_rdidx;
  assign regs_1_MPORT_4_mask = io_rdwmask_1;
  assign regs_1_MPORT_4_en = io_rdwen;
  assign regs_2_MPORT_en = 1'h1;
  assign regs_2_MPORT_addr = io_rs1idx;
  assign regs_2_MPORT_data = regs_2[regs_2_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_2_MPORT_1_en = 1'h1;
  assign regs_2_MPORT_1_addr = io_rs2idx;
  assign regs_2_MPORT_1_data = regs_2[regs_2_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_2_MPORT_2_en = 1'h1;
  assign regs_2_MPORT_2_addr = io_rs3idx;
  assign regs_2_MPORT_2_data = regs_2[regs_2_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_2_MPORT_3_en = 1'h1;
  assign regs_2_MPORT_3_addr = 5'h0;
  assign regs_2_MPORT_3_data = regs_2[regs_2_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_2_MPORT_4_data = io_rd_2;
  assign regs_2_MPORT_4_addr = io_rdidx;
  assign regs_2_MPORT_4_mask = io_rdwmask_2;
  assign regs_2_MPORT_4_en = io_rdwen;
  assign regs_3_MPORT_en = 1'h1;
  assign regs_3_MPORT_addr = io_rs1idx;
  assign regs_3_MPORT_data = regs_3[regs_3_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_3_MPORT_1_en = 1'h1;
  assign regs_3_MPORT_1_addr = io_rs2idx;
  assign regs_3_MPORT_1_data = regs_3[regs_3_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_3_MPORT_2_en = 1'h1;
  assign regs_3_MPORT_2_addr = io_rs3idx;
  assign regs_3_MPORT_2_data = regs_3[regs_3_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_3_MPORT_3_en = 1'h1;
  assign regs_3_MPORT_3_addr = 5'h0;
  assign regs_3_MPORT_3_data = regs_3[regs_3_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_3_MPORT_4_data = io_rd_3;
  assign regs_3_MPORT_4_addr = io_rdidx;
  assign regs_3_MPORT_4_mask = io_rdwmask_3;
  assign regs_3_MPORT_4_en = io_rdwen;
  assign regs_4_MPORT_en = 1'h1;
  assign regs_4_MPORT_addr = io_rs1idx;
  assign regs_4_MPORT_data = regs_4[regs_4_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_4_MPORT_1_en = 1'h1;
  assign regs_4_MPORT_1_addr = io_rs2idx;
  assign regs_4_MPORT_1_data = regs_4[regs_4_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_4_MPORT_2_en = 1'h1;
  assign regs_4_MPORT_2_addr = io_rs3idx;
  assign regs_4_MPORT_2_data = regs_4[regs_4_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_4_MPORT_3_en = 1'h1;
  assign regs_4_MPORT_3_addr = 5'h0;
  assign regs_4_MPORT_3_data = regs_4[regs_4_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_4_MPORT_4_data = io_rd_4;
  assign regs_4_MPORT_4_addr = io_rdidx;
  assign regs_4_MPORT_4_mask = io_rdwmask_4;
  assign regs_4_MPORT_4_en = io_rdwen;
  assign regs_5_MPORT_en = 1'h1;
  assign regs_5_MPORT_addr = io_rs1idx;
  assign regs_5_MPORT_data = regs_5[regs_5_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_5_MPORT_1_en = 1'h1;
  assign regs_5_MPORT_1_addr = io_rs2idx;
  assign regs_5_MPORT_1_data = regs_5[regs_5_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_5_MPORT_2_en = 1'h1;
  assign regs_5_MPORT_2_addr = io_rs3idx;
  assign regs_5_MPORT_2_data = regs_5[regs_5_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_5_MPORT_3_en = 1'h1;
  assign regs_5_MPORT_3_addr = 5'h0;
  assign regs_5_MPORT_3_data = regs_5[regs_5_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_5_MPORT_4_data = io_rd_5;
  assign regs_5_MPORT_4_addr = io_rdidx;
  assign regs_5_MPORT_4_mask = io_rdwmask_5;
  assign regs_5_MPORT_4_en = io_rdwen;
  assign regs_6_MPORT_en = 1'h1;
  assign regs_6_MPORT_addr = io_rs1idx;
  assign regs_6_MPORT_data = regs_6[regs_6_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_6_MPORT_1_en = 1'h1;
  assign regs_6_MPORT_1_addr = io_rs2idx;
  assign regs_6_MPORT_1_data = regs_6[regs_6_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_6_MPORT_2_en = 1'h1;
  assign regs_6_MPORT_2_addr = io_rs3idx;
  assign regs_6_MPORT_2_data = regs_6[regs_6_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_6_MPORT_3_en = 1'h1;
  assign regs_6_MPORT_3_addr = 5'h0;
  assign regs_6_MPORT_3_data = regs_6[regs_6_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_6_MPORT_4_data = io_rd_6;
  assign regs_6_MPORT_4_addr = io_rdidx;
  assign regs_6_MPORT_4_mask = io_rdwmask_6;
  assign regs_6_MPORT_4_en = io_rdwen;
  assign regs_7_MPORT_en = 1'h1;
  assign regs_7_MPORT_addr = io_rs1idx;
  assign regs_7_MPORT_data = regs_7[regs_7_MPORT_addr]; // @[regfile.scala 49:17]
  assign regs_7_MPORT_1_en = 1'h1;
  assign regs_7_MPORT_1_addr = io_rs2idx;
  assign regs_7_MPORT_1_data = regs_7[regs_7_MPORT_1_addr]; // @[regfile.scala 49:17]
  assign regs_7_MPORT_2_en = 1'h1;
  assign regs_7_MPORT_2_addr = io_rs3idx;
  assign regs_7_MPORT_2_data = regs_7[regs_7_MPORT_2_addr]; // @[regfile.scala 49:17]
  assign regs_7_MPORT_3_en = 1'h1;
  assign regs_7_MPORT_3_addr = 5'h0;
  assign regs_7_MPORT_3_data = regs_7[regs_7_MPORT_3_addr]; // @[regfile.scala 49:17]
  assign regs_7_MPORT_4_data = io_rd_7;
  assign regs_7_MPORT_4_addr = io_rdidx;
  assign regs_7_MPORT_4_mask = io_rdwmask_7;
  assign regs_7_MPORT_4_en = io_rdwen;
  assign io_v0_0 = regs_0_MPORT_3_data; // @[regfile.scala 54:9]
  assign io_rs1_0 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_0 : regs_0_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_1 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_1 : regs_1_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_2 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_2 : regs_2_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_3 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_3 : regs_3_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_4 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_4 : regs_4_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_5 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_5 : regs_5_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_6 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_6 : regs_6_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs1_7 = io_rs1idx == io_rdidx & io_rdwen ? io_rd_7 : regs_7_MPORT_data; // @[regfile.scala 51:16]
  assign io_rs2_0 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_0 : regs_0_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_1 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_1 : regs_1_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_2 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_2 : regs_2_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_3 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_3 : regs_3_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_4 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_4 : regs_4_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_5 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_5 : regs_5_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_6 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_6 : regs_6_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs2_7 = io_rs2idx == io_rdidx & io_rdwen ? io_rd_7 : regs_7_MPORT_1_data; // @[regfile.scala 52:16]
  assign io_rs3_0 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_0 : regs_0_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_1 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_1 : regs_1_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_2 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_2 : regs_2_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_3 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_3 : regs_3_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_4 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_4 : regs_4_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_5 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_5 : regs_5_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_6 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_6 : regs_6_MPORT_2_data; // @[regfile.scala 53:16]
  assign io_rs3_7 = io_rs3idx == io_rdidx & io_rdwen ? io_rd_7 : regs_7_MPORT_2_data; // @[regfile.scala 53:16]
  always @(posedge clock) begin
    if (regs_0_MPORT_4_en & regs_0_MPORT_4_mask) begin
      regs_0[regs_0_MPORT_4_addr] <= regs_0_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_1_MPORT_4_en & regs_1_MPORT_4_mask) begin
      regs_1[regs_1_MPORT_4_addr] <= regs_1_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_2_MPORT_4_en & regs_2_MPORT_4_mask) begin
      regs_2[regs_2_MPORT_4_addr] <= regs_2_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_3_MPORT_4_en & regs_3_MPORT_4_mask) begin
      regs_3[regs_3_MPORT_4_addr] <= regs_3_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_4_MPORT_4_en & regs_4_MPORT_4_mask) begin
      regs_4[regs_4_MPORT_4_addr] <= regs_4_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_5_MPORT_4_en & regs_5_MPORT_4_mask) begin
      regs_5[regs_5_MPORT_4_addr] <= regs_5_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_6_MPORT_4_en & regs_6_MPORT_4_mask) begin
      regs_6[regs_6_MPORT_4_addr] <= regs_6_MPORT_4_data; // @[regfile.scala 49:17]
    end
    if (regs_7_MPORT_4_en & regs_7_MPORT_4_mask) begin
      regs_7[regs_7_MPORT_4_addr] <= regs_7_MPORT_4_data; // @[regfile.scala 49:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_0[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_1[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_2[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_3[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_4[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_5[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_6[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs_7[initvar] = _RAND_7[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile(
  input         clock,
  output [31:0] io_rs1,
  output [31:0] io_rs2,
  output [31:0] io_rs3,
  input  [4:0]  io_rs1idx,
  input  [4:0]  io_rs2idx,
  input  [4:0]  io_rs3idx,
  input  [31:0] io_rd,
  input  [4:0]  io_rdidx,
  input         io_rdwen
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] regs [0:31]; // @[regfile.scala 23:17]
  wire  regs_io_rs1_MPORT_en; // @[regfile.scala 23:17]
  wire [4:0] regs_io_rs1_MPORT_addr; // @[regfile.scala 23:17]
  wire [31:0] regs_io_rs1_MPORT_data; // @[regfile.scala 23:17]
  wire  regs_io_rs2_MPORT_en; // @[regfile.scala 23:17]
  wire [4:0] regs_io_rs2_MPORT_addr; // @[regfile.scala 23:17]
  wire [31:0] regs_io_rs2_MPORT_data; // @[regfile.scala 23:17]
  wire  regs_io_rs3_MPORT_en; // @[regfile.scala 23:17]
  wire [4:0] regs_io_rs3_MPORT_addr; // @[regfile.scala 23:17]
  wire [31:0] regs_io_rs3_MPORT_data; // @[regfile.scala 23:17]
  wire  regs_io_x1_MPORT_en; // @[regfile.scala 23:17]
  wire [4:0] regs_io_x1_MPORT_addr; // @[regfile.scala 23:17]
  wire [31:0] regs_io_x1_MPORT_data; // @[regfile.scala 23:17]
  wire [31:0] regs_MPORT_data; // @[regfile.scala 23:17]
  wire [4:0] regs_MPORT_addr; // @[regfile.scala 23:17]
  wire  regs_MPORT_mask; // @[regfile.scala 23:17]
  wire  regs_MPORT_en; // @[regfile.scala 23:17]
  wire [31:0] _io_rs1_T_3 = |io_rs1idx ? regs_io_rs1_MPORT_data : 32'h0; // @[regfile.scala 24:60]
  wire [31:0] _io_rs2_T_3 = |io_rs2idx ? regs_io_rs2_MPORT_data : 32'h0; // @[regfile.scala 25:60]
  wire [31:0] _io_rs3_T_3 = |io_rs3idx ? regs_io_rs3_MPORT_data : 32'h0; // @[regfile.scala 26:60]
  wire  _T = |io_rdidx; // @[regfile.scala 28:29]
  assign regs_io_rs1_MPORT_en = 1'h1;
  assign regs_io_rs1_MPORT_addr = io_rs1idx;
  assign regs_io_rs1_MPORT_data = regs[regs_io_rs1_MPORT_addr]; // @[regfile.scala 23:17]
  assign regs_io_rs2_MPORT_en = 1'h1;
  assign regs_io_rs2_MPORT_addr = io_rs2idx;
  assign regs_io_rs2_MPORT_data = regs[regs_io_rs2_MPORT_addr]; // @[regfile.scala 23:17]
  assign regs_io_rs3_MPORT_en = 1'h1;
  assign regs_io_rs3_MPORT_addr = io_rs3idx;
  assign regs_io_rs3_MPORT_data = regs[regs_io_rs3_MPORT_addr]; // @[regfile.scala 23:17]
  assign regs_io_x1_MPORT_en = 1'h1;
  assign regs_io_x1_MPORT_addr = 5'h1;
  assign regs_io_x1_MPORT_data = regs[regs_io_x1_MPORT_addr]; // @[regfile.scala 23:17]
  assign regs_MPORT_data = io_rd;
  assign regs_MPORT_addr = io_rdidx;
  assign regs_MPORT_mask = 1'h1;
  assign regs_MPORT_en = io_rdwen & _T;
  assign io_rs1 = io_rs1idx == io_rdidx & io_rdwen ? io_rd : _io_rs1_T_3; // @[regfile.scala 24:16]
  assign io_rs2 = io_rs2idx == io_rdidx & io_rdwen ? io_rd : _io_rs2_T_3; // @[regfile.scala 25:16]
  assign io_rs3 = io_rs3idx == io_rdidx & io_rdwen ? io_rd : _io_rs3_T_3; // @[regfile.scala 26:16]
  always @(posedge clock) begin
    if (regs_MPORT_en & regs_MPORT_mask) begin
      regs[regs_MPORT_addr] <= regs_MPORT_data; // @[regfile.scala 23:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ImmGen(
  input  [31:0] io_inst,
  input  [2:0]  io_sel,
  output [31:0] io_out
);
  wire [11:0] Iimm = io_inst[31:20]; // @[regfile.scala 72:30]
  wire [11:0] Simm = {io_inst[31:25],io_inst[11:7]}; // @[regfile.scala 73:51]
  wire [12:0] Bimm = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[regfile.scala 74:86]
  wire [31:0] Uimm = {io_inst[31:12],12'h0}; // @[regfile.scala 75:46]
  wire [20:0] Jimm = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[regfile.scala 76:88]
  wire [31:0] Zimm = {27'h0,io_inst[19:15]}; // @[regfile.scala 77:45]
  wire [4:0] Imm2 = io_inst[24:20]; // @[regfile.scala 78:29]
  wire [4:0] Vimm = io_inst[19:15]; // @[regfile.scala 79:29]
  wire [20:0] _out_T_3 = 3'h5 == io_sel ? $signed(Jimm) : $signed({{9{Iimm[11]}},Iimm}); // @[Mux.scala 81:58]
  wire [20:0] _out_T_5 = 3'h1 == io_sel ? $signed({{9{Simm[11]}},Simm}) : $signed(_out_T_3); // @[Mux.scala 81:58]
  wire [20:0] _out_T_7 = 3'h2 == io_sel ? $signed({{8{Bimm[12]}},Bimm}) : $signed(_out_T_5); // @[Mux.scala 81:58]
  wire [31:0] _out_T_9 = 3'h3 == io_sel ? $signed(Uimm) : $signed({{11{_out_T_7[20]}},_out_T_7}); // @[Mux.scala 81:58]
  wire [31:0] _out_T_11 = 3'h4 == io_sel ? $signed({{27{Imm2[4]}},Imm2}) : $signed(_out_T_9); // @[Mux.scala 81:58]
  wire [31:0] _out_T_13 = 3'h7 == io_sel ? $signed(Zimm) : $signed(_out_T_11); // @[Mux.scala 81:58]
  assign io_out = 3'h6 == io_sel ? $signed({{27{Vimm[4]}},Vimm}) : $signed(_out_T_13); // @[regfile.scala 84:15]
endmodule
module operandCollector(
  input         clock,
  input  [31:0] io_control_inst,
  input  [1:0]  io_control_wid,
  input  [1:0]  io_control_branch,
  input  [1:0]  io_control_sel_alu2,
  input  [1:0]  io_control_sel_alu1,
  input         io_control_isvec,
  input  [1:0]  io_control_sel_alu3,
  input         io_control_mask,
  input  [2:0]  io_control_sel_imm,
  input  [4:0]  io_control_reg_idx1,
  input  [4:0]  io_control_reg_idx2,
  input  [4:0]  io_control_reg_idx3,
  input  [31:0] io_control_pc,
  output [31:0] io_alu_src1_0,
  output [31:0] io_alu_src1_1,
  output [31:0] io_alu_src1_2,
  output [31:0] io_alu_src1_3,
  output [31:0] io_alu_src1_4,
  output [31:0] io_alu_src1_5,
  output [31:0] io_alu_src1_6,
  output [31:0] io_alu_src1_7,
  output [31:0] io_alu_src2_0,
  output [31:0] io_alu_src2_1,
  output [31:0] io_alu_src2_2,
  output [31:0] io_alu_src2_3,
  output [31:0] io_alu_src2_4,
  output [31:0] io_alu_src2_5,
  output [31:0] io_alu_src2_6,
  output [31:0] io_alu_src2_7,
  output [31:0] io_alu_src3_0,
  output [31:0] io_alu_src3_1,
  output [31:0] io_alu_src3_2,
  output [31:0] io_alu_src3_3,
  output [31:0] io_alu_src3_4,
  output [31:0] io_alu_src3_5,
  output [31:0] io_alu_src3_6,
  output [31:0] io_alu_src3_7,
  output        io_mask_0,
  output        io_mask_1,
  output        io_mask_2,
  output        io_mask_3,
  output        io_mask_4,
  output        io_mask_5,
  output        io_mask_6,
  output        io_mask_7,
  input         io_writeScalarCtrl_valid,
  input  [31:0] io_writeScalarCtrl_bits_wb_wxd_rd,
  input         io_writeScalarCtrl_bits_wxd,
  input  [4:0]  io_writeScalarCtrl_bits_reg_idxw,
  input  [1:0]  io_writeScalarCtrl_bits_warp_id,
  input         io_writeVecCtrl_valid,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_0,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_1,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_2,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_3,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_4,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_5,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_6,
  input  [31:0] io_writeVecCtrl_bits_wb_wfd_rd_7,
  input         io_writeVecCtrl_bits_wfd_mask_0,
  input         io_writeVecCtrl_bits_wfd_mask_1,
  input         io_writeVecCtrl_bits_wfd_mask_2,
  input         io_writeVecCtrl_bits_wfd_mask_3,
  input         io_writeVecCtrl_bits_wfd_mask_4,
  input         io_writeVecCtrl_bits_wfd_mask_5,
  input         io_writeVecCtrl_bits_wfd_mask_6,
  input         io_writeVecCtrl_bits_wfd_mask_7,
  input         io_writeVecCtrl_bits_wfd,
  input  [4:0]  io_writeVecCtrl_bits_reg_idxw,
  input  [1:0]  io_writeVecCtrl_bits_warp_id
);
  wire  FloatRegFile_clock; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_v0_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs1_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs2_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rs3_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_io_rs1idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_io_rs2idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_io_rs3idx; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_io_rd_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_io_rdidx; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwen; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_0; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_1; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_2; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_3; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_4; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_5; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_6; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_io_rdwmask_7; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_clock; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_v0_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs1_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs2_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rs3_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_1_io_rs1idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_1_io_rs2idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_1_io_rs3idx; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_1_io_rd_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_1_io_rdidx; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwen; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_0; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_1; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_2; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_3; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_4; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_5; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_6; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_1_io_rdwmask_7; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_clock; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_v0_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs1_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs2_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rs3_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_2_io_rs1idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_2_io_rs2idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_2_io_rs3idx; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_2_io_rd_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_2_io_rdidx; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwen; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_0; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_1; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_2; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_3; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_4; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_5; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_6; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_2_io_rdwmask_7; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_clock; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_v0_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs1_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs2_7; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rs3_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_3_io_rs1idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_3_io_rs2idx; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_3_io_rs3idx; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_0; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_1; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_2; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_3; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_4; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_5; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_6; // @[operandCollector.scala 34:54]
  wire [31:0] FloatRegFile_3_io_rd_7; // @[operandCollector.scala 34:54]
  wire [4:0] FloatRegFile_3_io_rdidx; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwen; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_0; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_1; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_2; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_3; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_4; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_5; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_6; // @[operandCollector.scala 34:54]
  wire  FloatRegFile_3_io_rdwmask_7; // @[operandCollector.scala 34:54]
  wire  RegFile_clock; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_io_rs1; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_io_rs2; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_io_rs3; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_io_rs1idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_io_rs2idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_io_rs3idx; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_io_rd; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_io_rdidx; // @[operandCollector.scala 35:54]
  wire  RegFile_io_rdwen; // @[operandCollector.scala 35:54]
  wire  RegFile_1_clock; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_1_io_rs1; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_1_io_rs2; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_1_io_rs3; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_1_io_rs1idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_1_io_rs2idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_1_io_rs3idx; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_1_io_rd; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_1_io_rdidx; // @[operandCollector.scala 35:54]
  wire  RegFile_1_io_rdwen; // @[operandCollector.scala 35:54]
  wire  RegFile_2_clock; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_2_io_rs1; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_2_io_rs2; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_2_io_rs3; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_2_io_rs1idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_2_io_rs2idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_2_io_rs3idx; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_2_io_rd; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_2_io_rdidx; // @[operandCollector.scala 35:54]
  wire  RegFile_2_io_rdwen; // @[operandCollector.scala 35:54]
  wire  RegFile_3_clock; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_3_io_rs1; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_3_io_rs2; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_3_io_rs3; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_3_io_rs1idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_3_io_rs2idx; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_3_io_rs3idx; // @[operandCollector.scala 35:54]
  wire [31:0] RegFile_3_io_rd; // @[operandCollector.scala 35:54]
  wire [4:0] RegFile_3_io_rdidx; // @[operandCollector.scala 35:54]
  wire  RegFile_3_io_rdwen; // @[operandCollector.scala 35:54]
  wire [31:0] imm_io_inst; // @[operandCollector.scala 36:17]
  wire [2:0] imm_io_sel; // @[operandCollector.scala 36:17]
  wire [31:0] imm_io_out; // @[operandCollector.scala 36:17]
  wire [31:0] vectorRegFile_0_rs1_0 = FloatRegFile_io_rs1_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_0 = FloatRegFile_1_io_rs1_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_9 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_0 : vectorRegFile_0_rs1_0; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_0 = FloatRegFile_2_io_rs1_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_10 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_0 : _GEN_9; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_0 = FloatRegFile_3_io_rs1_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_11 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_0 : _GEN_10; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_0_rs1 = RegFile_io_rs1; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] scalarRegFile_1_rs1 = RegFile_1_io_rs1; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_13 = 2'h1 == io_control_wid ? scalarRegFile_1_rs1 : scalarRegFile_0_rs1; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_2_rs1 = RegFile_2_io_rs1; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_14 = 2'h2 == io_control_wid ? scalarRegFile_2_rs1 : _GEN_13; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_3_rs1 = RegFile_3_io_rs1; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_15 = 2'h3 == io_control_wid ? scalarRegFile_3_rs1 : _GEN_14; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_0_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_11 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_0_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] scalarRegFile_0_rs2 = RegFile_io_rs2; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] scalarRegFile_1_rs2 = RegFile_1_io_rs2; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_17 = 2'h1 == io_control_wid ? scalarRegFile_1_rs2 : scalarRegFile_0_rs2; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_2_rs2 = RegFile_2_io_rs2; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_18 = 2'h2 == io_control_wid ? scalarRegFile_2_rs2 : _GEN_17; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_3_rs2 = RegFile_3_io_rs2; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_19 = 2'h3 == io_control_wid ? scalarRegFile_3_rs2 : _GEN_18; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_0_T_1 = 2'h3 == io_control_sel_alu2 ? imm_io_out : _GEN_19; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_0 = FloatRegFile_io_rs2_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_0 = FloatRegFile_1_io_rs2_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_21 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_0 : vectorRegFile_0_rs2_0; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_0 = FloatRegFile_2_io_rs2_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_22 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_0 : _GEN_21; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_0 = FloatRegFile_3_io_rs2_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_23 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_0 : _GEN_22; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_0_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_23 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_0_T_2 = imm_io_out + _GEN_15; // @[operandCollector.scala 67:107]
  wire [31:0] _io_alu_src3_0_T_4 = io_control_pc + imm_io_out; // @[operandCollector.scala 67:157]
  wire [31:0] _io_alu_src3_0_T_5 = io_control_branch == 2'h3 ? _io_alu_src3_0_T_2 : _io_alu_src3_0_T_4; // @[operandCollector.scala 67:71]
  wire [31:0] vectorRegFile_0_rs3_0 = FloatRegFile_io_rs3_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_0 = FloatRegFile_1_io_rs3_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_25 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_0 : vectorRegFile_0_rs3_0; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_0 = FloatRegFile_2_io_rs3_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_26 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_0 : _GEN_25; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_0 = FloatRegFile_3_io_rs3_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_27 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_0 : _GEN_26; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_0_T_6 = io_control_isvec ? _GEN_27 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_0_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_27 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_0_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_0_T_6 : _io_alu_src3_0_T_8; // @[Mux.scala 81:58]
  wire [31:0] scalarRegFile_0_rs3 = RegFile_io_rs3; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] scalarRegFile_1_rs3 = RegFile_1_io_rs3; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_29 = 2'h1 == io_control_wid ? scalarRegFile_1_rs3 : scalarRegFile_0_rs3; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_2_rs3 = RegFile_2_io_rs3; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_30 = 2'h2 == io_control_wid ? scalarRegFile_2_rs3 : _GEN_29; // @[Mux.scala 81:{58,58}]
  wire [31:0] scalarRegFile_3_rs3 = RegFile_3_io_rs3; // @[operandCollector.scala 35:{28,28}]
  wire [31:0] _GEN_31 = 2'h3 == io_control_wid ? scalarRegFile_3_rs3 : _GEN_30; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_0_v0_0 = FloatRegFile_io_v0_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_v0_0 = FloatRegFile_1_io_v0_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_33 = 2'h1 == io_control_wid ? vectorRegFile_1_v0_0 : vectorRegFile_0_v0_0; // @[operandCollector.scala 68:{78,78}]
  wire [31:0] vectorRegFile_2_v0_0 = FloatRegFile_2_io_v0_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_34 = 2'h2 == io_control_wid ? vectorRegFile_2_v0_0 : _GEN_33; // @[operandCollector.scala 68:{78,78}]
  wire [31:0] vectorRegFile_3_v0_0 = FloatRegFile_3_io_v0_0; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_35 = 2'h3 == io_control_wid ? vectorRegFile_3_v0_0 : _GEN_34; // @[operandCollector.scala 68:{78,78}]
  wire [31:0] vectorRegFile_0_rs1_1 = FloatRegFile_io_rs1_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_1 = FloatRegFile_1_io_rs1_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_37 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_1 : vectorRegFile_0_rs1_1; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_1 = FloatRegFile_2_io_rs1_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_38 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_1 : _GEN_37; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_1 = FloatRegFile_3_io_rs1_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_39 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_1 : _GEN_38; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_1_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_39 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_1_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_1_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_1 = FloatRegFile_io_rs2_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_1 = FloatRegFile_1_io_rs2_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_41 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_1 : vectorRegFile_0_rs2_1; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_1 = FloatRegFile_2_io_rs2_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_42 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_1 : _GEN_41; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_1 = FloatRegFile_3_io_rs2_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_43 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_1 : _GEN_42; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_1_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_43 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_1 = FloatRegFile_io_rs3_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_1 = FloatRegFile_1_io_rs3_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_45 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_1 : vectorRegFile_0_rs3_1; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_1 = FloatRegFile_2_io_rs3_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_46 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_1 : _GEN_45; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_1 = FloatRegFile_3_io_rs3_1; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_47 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_1 : _GEN_46; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_1_T_6 = io_control_isvec ? _GEN_47 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_1_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_47 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_1_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_1_T_6 : _io_alu_src3_1_T_8; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs1_2 = FloatRegFile_io_rs1_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_2 = FloatRegFile_1_io_rs1_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_49 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_2 : vectorRegFile_0_rs1_2; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_2 = FloatRegFile_2_io_rs1_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_50 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_2 : _GEN_49; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_2 = FloatRegFile_3_io_rs1_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_51 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_2 : _GEN_50; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_2_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_51 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_2_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_2_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_2 = FloatRegFile_io_rs2_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_2 = FloatRegFile_1_io_rs2_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_53 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_2 : vectorRegFile_0_rs2_2; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_2 = FloatRegFile_2_io_rs2_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_54 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_2 : _GEN_53; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_2 = FloatRegFile_3_io_rs2_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_55 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_2 : _GEN_54; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_2_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_55 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_2 = FloatRegFile_io_rs3_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_2 = FloatRegFile_1_io_rs3_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_57 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_2 : vectorRegFile_0_rs3_2; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_2 = FloatRegFile_2_io_rs3_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_58 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_2 : _GEN_57; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_2 = FloatRegFile_3_io_rs3_2; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_59 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_2 : _GEN_58; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_2_T_6 = io_control_isvec ? _GEN_59 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_2_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_59 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_2_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_2_T_6 : _io_alu_src3_2_T_8; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs1_3 = FloatRegFile_io_rs1_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_3 = FloatRegFile_1_io_rs1_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_61 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_3 : vectorRegFile_0_rs1_3; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_3 = FloatRegFile_2_io_rs1_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_62 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_3 : _GEN_61; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_3 = FloatRegFile_3_io_rs1_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_63 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_3 : _GEN_62; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_3_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_63 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_3_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_3_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_3 = FloatRegFile_io_rs2_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_3 = FloatRegFile_1_io_rs2_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_65 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_3 : vectorRegFile_0_rs2_3; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_3 = FloatRegFile_2_io_rs2_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_66 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_3 : _GEN_65; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_3 = FloatRegFile_3_io_rs2_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_67 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_3 : _GEN_66; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_3_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_67 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_3 = FloatRegFile_io_rs3_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_3 = FloatRegFile_1_io_rs3_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_69 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_3 : vectorRegFile_0_rs3_3; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_3 = FloatRegFile_2_io_rs3_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_70 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_3 : _GEN_69; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_3 = FloatRegFile_3_io_rs3_3; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_71 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_3 : _GEN_70; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_3_T_6 = io_control_isvec ? _GEN_71 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_3_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_71 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_3_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_3_T_6 : _io_alu_src3_3_T_8; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs1_4 = FloatRegFile_io_rs1_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_4 = FloatRegFile_1_io_rs1_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_73 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_4 : vectorRegFile_0_rs1_4; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_4 = FloatRegFile_2_io_rs1_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_74 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_4 : _GEN_73; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_4 = FloatRegFile_3_io_rs1_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_75 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_4 : _GEN_74; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_4_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_75 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_4_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_4_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_4 = FloatRegFile_io_rs2_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_4 = FloatRegFile_1_io_rs2_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_77 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_4 : vectorRegFile_0_rs2_4; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_4 = FloatRegFile_2_io_rs2_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_78 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_4 : _GEN_77; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_4 = FloatRegFile_3_io_rs2_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_79 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_4 : _GEN_78; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_4_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_79 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_4 = FloatRegFile_io_rs3_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_4 = FloatRegFile_1_io_rs3_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_81 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_4 : vectorRegFile_0_rs3_4; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_4 = FloatRegFile_2_io_rs3_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_82 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_4 : _GEN_81; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_4 = FloatRegFile_3_io_rs3_4; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_83 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_4 : _GEN_82; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_4_T_6 = io_control_isvec ? _GEN_83 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_4_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_83 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_4_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_4_T_6 : _io_alu_src3_4_T_8; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs1_5 = FloatRegFile_io_rs1_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_5 = FloatRegFile_1_io_rs1_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_85 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_5 : vectorRegFile_0_rs1_5; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_5 = FloatRegFile_2_io_rs1_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_86 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_5 : _GEN_85; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_5 = FloatRegFile_3_io_rs1_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_87 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_5 : _GEN_86; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_5_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_87 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_5_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_5_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_5 = FloatRegFile_io_rs2_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_5 = FloatRegFile_1_io_rs2_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_89 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_5 : vectorRegFile_0_rs2_5; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_5 = FloatRegFile_2_io_rs2_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_90 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_5 : _GEN_89; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_5 = FloatRegFile_3_io_rs2_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_91 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_5 : _GEN_90; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_5_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_91 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_5 = FloatRegFile_io_rs3_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_5 = FloatRegFile_1_io_rs3_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_93 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_5 : vectorRegFile_0_rs3_5; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_5 = FloatRegFile_2_io_rs3_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_94 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_5 : _GEN_93; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_5 = FloatRegFile_3_io_rs3_5; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_95 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_5 : _GEN_94; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_5_T_6 = io_control_isvec ? _GEN_95 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_5_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_95 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_5_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_5_T_6 : _io_alu_src3_5_T_8; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs1_6 = FloatRegFile_io_rs1_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_6 = FloatRegFile_1_io_rs1_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_97 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_6 : vectorRegFile_0_rs1_6; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_6 = FloatRegFile_2_io_rs1_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_98 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_6 : _GEN_97; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_6 = FloatRegFile_3_io_rs1_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_99 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_6 : _GEN_98; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_6_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_99 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_6_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_6_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_6 = FloatRegFile_io_rs2_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_6 = FloatRegFile_1_io_rs2_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_101 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_6 : vectorRegFile_0_rs2_6; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_6 = FloatRegFile_2_io_rs2_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_102 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_6 : _GEN_101; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_6 = FloatRegFile_3_io_rs2_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_103 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_6 : _GEN_102; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_6_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_103 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_6 = FloatRegFile_io_rs3_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_6 = FloatRegFile_1_io_rs3_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_105 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_6 : vectorRegFile_0_rs3_6; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_6 = FloatRegFile_2_io_rs3_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_106 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_6 : _GEN_105; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_6 = FloatRegFile_3_io_rs3_6; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_107 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_6 : _GEN_106; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_6_T_6 = io_control_isvec ? _GEN_107 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_6_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_107 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_6_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_6_T_6 : _io_alu_src3_6_T_8; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs1_7 = FloatRegFile_io_rs1_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs1_7 = FloatRegFile_1_io_rs1_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_109 = 2'h1 == io_control_wid ? vectorRegFile_1_rs1_7 : vectorRegFile_0_rs1_7; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs1_7 = FloatRegFile_2_io_rs1_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_110 = 2'h2 == io_control_wid ? vectorRegFile_2_rs1_7 : _GEN_109; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs1_7 = FloatRegFile_3_io_rs1_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_111 = 2'h3 == io_control_wid ? vectorRegFile_3_rs1_7 : _GEN_110; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src1_7_T_1 = 2'h2 == io_control_sel_alu1 ? _GEN_111 : _GEN_15; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src1_7_T_3 = 2'h3 == io_control_sel_alu1 ? imm_io_out : _io_alu_src1_7_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs2_7 = FloatRegFile_io_rs2_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs2_7 = FloatRegFile_1_io_rs2_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_113 = 2'h1 == io_control_wid ? vectorRegFile_1_rs2_7 : vectorRegFile_0_rs2_7; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_2_rs2_7 = FloatRegFile_2_io_rs2_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_114 = 2'h2 == io_control_wid ? vectorRegFile_2_rs2_7 : _GEN_113; // @[Mux.scala 81:{58,58}]
  wire [31:0] vectorRegFile_3_rs2_7 = FloatRegFile_3_io_rs2_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_115 = 2'h3 == io_control_wid ? vectorRegFile_3_rs2_7 : _GEN_114; // @[Mux.scala 81:{58,58}]
  wire [31:0] _io_alu_src2_7_T_3 = 2'h2 == io_control_sel_alu2 ? _GEN_115 : _io_alu_src2_0_T_1; // @[Mux.scala 81:58]
  wire [31:0] vectorRegFile_0_rs3_7 = FloatRegFile_io_rs3_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] vectorRegFile_1_rs3_7 = FloatRegFile_1_io_rs3_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_117 = 2'h1 == io_control_wid ? vectorRegFile_1_rs3_7 : vectorRegFile_0_rs3_7; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_2_rs3_7 = FloatRegFile_2_io_rs3_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_118 = 2'h2 == io_control_wid ? vectorRegFile_2_rs3_7 : _GEN_117; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] vectorRegFile_3_rs3_7 = FloatRegFile_3_io_rs3_7; // @[operandCollector.scala 34:{28,28}]
  wire [31:0] _GEN_119 = 2'h3 == io_control_wid ? vectorRegFile_3_rs3_7 : _GEN_118; // @[operandCollector.scala 67:{227,227}]
  wire [31:0] _io_alu_src3_7_T_6 = io_control_isvec ? _GEN_119 : _GEN_19; // @[operandCollector.scala 67:227]
  wire [31:0] _io_alu_src3_7_T_8 = 2'h1 == io_control_sel_alu3 ? _GEN_119 : _io_alu_src3_0_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_alu_src3_7_T_10 = 2'h3 == io_control_sel_alu3 ? _io_alu_src3_7_T_6 : _io_alu_src3_7_T_8; // @[Mux.scala 81:58]
  FloatRegFile FloatRegFile ( // @[operandCollector.scala 34:54]
    .clock(FloatRegFile_clock),
    .io_v0_0(FloatRegFile_io_v0_0),
    .io_rs1_0(FloatRegFile_io_rs1_0),
    .io_rs1_1(FloatRegFile_io_rs1_1),
    .io_rs1_2(FloatRegFile_io_rs1_2),
    .io_rs1_3(FloatRegFile_io_rs1_3),
    .io_rs1_4(FloatRegFile_io_rs1_4),
    .io_rs1_5(FloatRegFile_io_rs1_5),
    .io_rs1_6(FloatRegFile_io_rs1_6),
    .io_rs1_7(FloatRegFile_io_rs1_7),
    .io_rs2_0(FloatRegFile_io_rs2_0),
    .io_rs2_1(FloatRegFile_io_rs2_1),
    .io_rs2_2(FloatRegFile_io_rs2_2),
    .io_rs2_3(FloatRegFile_io_rs2_3),
    .io_rs2_4(FloatRegFile_io_rs2_4),
    .io_rs2_5(FloatRegFile_io_rs2_5),
    .io_rs2_6(FloatRegFile_io_rs2_6),
    .io_rs2_7(FloatRegFile_io_rs2_7),
    .io_rs3_0(FloatRegFile_io_rs3_0),
    .io_rs3_1(FloatRegFile_io_rs3_1),
    .io_rs3_2(FloatRegFile_io_rs3_2),
    .io_rs3_3(FloatRegFile_io_rs3_3),
    .io_rs3_4(FloatRegFile_io_rs3_4),
    .io_rs3_5(FloatRegFile_io_rs3_5),
    .io_rs3_6(FloatRegFile_io_rs3_6),
    .io_rs3_7(FloatRegFile_io_rs3_7),
    .io_rs1idx(FloatRegFile_io_rs1idx),
    .io_rs2idx(FloatRegFile_io_rs2idx),
    .io_rs3idx(FloatRegFile_io_rs3idx),
    .io_rd_0(FloatRegFile_io_rd_0),
    .io_rd_1(FloatRegFile_io_rd_1),
    .io_rd_2(FloatRegFile_io_rd_2),
    .io_rd_3(FloatRegFile_io_rd_3),
    .io_rd_4(FloatRegFile_io_rd_4),
    .io_rd_5(FloatRegFile_io_rd_5),
    .io_rd_6(FloatRegFile_io_rd_6),
    .io_rd_7(FloatRegFile_io_rd_7),
    .io_rdidx(FloatRegFile_io_rdidx),
    .io_rdwen(FloatRegFile_io_rdwen),
    .io_rdwmask_0(FloatRegFile_io_rdwmask_0),
    .io_rdwmask_1(FloatRegFile_io_rdwmask_1),
    .io_rdwmask_2(FloatRegFile_io_rdwmask_2),
    .io_rdwmask_3(FloatRegFile_io_rdwmask_3),
    .io_rdwmask_4(FloatRegFile_io_rdwmask_4),
    .io_rdwmask_5(FloatRegFile_io_rdwmask_5),
    .io_rdwmask_6(FloatRegFile_io_rdwmask_6),
    .io_rdwmask_7(FloatRegFile_io_rdwmask_7)
  );
  FloatRegFile FloatRegFile_1 ( // @[operandCollector.scala 34:54]
    .clock(FloatRegFile_1_clock),
    .io_v0_0(FloatRegFile_1_io_v0_0),
    .io_rs1_0(FloatRegFile_1_io_rs1_0),
    .io_rs1_1(FloatRegFile_1_io_rs1_1),
    .io_rs1_2(FloatRegFile_1_io_rs1_2),
    .io_rs1_3(FloatRegFile_1_io_rs1_3),
    .io_rs1_4(FloatRegFile_1_io_rs1_4),
    .io_rs1_5(FloatRegFile_1_io_rs1_5),
    .io_rs1_6(FloatRegFile_1_io_rs1_6),
    .io_rs1_7(FloatRegFile_1_io_rs1_7),
    .io_rs2_0(FloatRegFile_1_io_rs2_0),
    .io_rs2_1(FloatRegFile_1_io_rs2_1),
    .io_rs2_2(FloatRegFile_1_io_rs2_2),
    .io_rs2_3(FloatRegFile_1_io_rs2_3),
    .io_rs2_4(FloatRegFile_1_io_rs2_4),
    .io_rs2_5(FloatRegFile_1_io_rs2_5),
    .io_rs2_6(FloatRegFile_1_io_rs2_6),
    .io_rs2_7(FloatRegFile_1_io_rs2_7),
    .io_rs3_0(FloatRegFile_1_io_rs3_0),
    .io_rs3_1(FloatRegFile_1_io_rs3_1),
    .io_rs3_2(FloatRegFile_1_io_rs3_2),
    .io_rs3_3(FloatRegFile_1_io_rs3_3),
    .io_rs3_4(FloatRegFile_1_io_rs3_4),
    .io_rs3_5(FloatRegFile_1_io_rs3_5),
    .io_rs3_6(FloatRegFile_1_io_rs3_6),
    .io_rs3_7(FloatRegFile_1_io_rs3_7),
    .io_rs1idx(FloatRegFile_1_io_rs1idx),
    .io_rs2idx(FloatRegFile_1_io_rs2idx),
    .io_rs3idx(FloatRegFile_1_io_rs3idx),
    .io_rd_0(FloatRegFile_1_io_rd_0),
    .io_rd_1(FloatRegFile_1_io_rd_1),
    .io_rd_2(FloatRegFile_1_io_rd_2),
    .io_rd_3(FloatRegFile_1_io_rd_3),
    .io_rd_4(FloatRegFile_1_io_rd_4),
    .io_rd_5(FloatRegFile_1_io_rd_5),
    .io_rd_6(FloatRegFile_1_io_rd_6),
    .io_rd_7(FloatRegFile_1_io_rd_7),
    .io_rdidx(FloatRegFile_1_io_rdidx),
    .io_rdwen(FloatRegFile_1_io_rdwen),
    .io_rdwmask_0(FloatRegFile_1_io_rdwmask_0),
    .io_rdwmask_1(FloatRegFile_1_io_rdwmask_1),
    .io_rdwmask_2(FloatRegFile_1_io_rdwmask_2),
    .io_rdwmask_3(FloatRegFile_1_io_rdwmask_3),
    .io_rdwmask_4(FloatRegFile_1_io_rdwmask_4),
    .io_rdwmask_5(FloatRegFile_1_io_rdwmask_5),
    .io_rdwmask_6(FloatRegFile_1_io_rdwmask_6),
    .io_rdwmask_7(FloatRegFile_1_io_rdwmask_7)
  );
  FloatRegFile FloatRegFile_2 ( // @[operandCollector.scala 34:54]
    .clock(FloatRegFile_2_clock),
    .io_v0_0(FloatRegFile_2_io_v0_0),
    .io_rs1_0(FloatRegFile_2_io_rs1_0),
    .io_rs1_1(FloatRegFile_2_io_rs1_1),
    .io_rs1_2(FloatRegFile_2_io_rs1_2),
    .io_rs1_3(FloatRegFile_2_io_rs1_3),
    .io_rs1_4(FloatRegFile_2_io_rs1_4),
    .io_rs1_5(FloatRegFile_2_io_rs1_5),
    .io_rs1_6(FloatRegFile_2_io_rs1_6),
    .io_rs1_7(FloatRegFile_2_io_rs1_7),
    .io_rs2_0(FloatRegFile_2_io_rs2_0),
    .io_rs2_1(FloatRegFile_2_io_rs2_1),
    .io_rs2_2(FloatRegFile_2_io_rs2_2),
    .io_rs2_3(FloatRegFile_2_io_rs2_3),
    .io_rs2_4(FloatRegFile_2_io_rs2_4),
    .io_rs2_5(FloatRegFile_2_io_rs2_5),
    .io_rs2_6(FloatRegFile_2_io_rs2_6),
    .io_rs2_7(FloatRegFile_2_io_rs2_7),
    .io_rs3_0(FloatRegFile_2_io_rs3_0),
    .io_rs3_1(FloatRegFile_2_io_rs3_1),
    .io_rs3_2(FloatRegFile_2_io_rs3_2),
    .io_rs3_3(FloatRegFile_2_io_rs3_3),
    .io_rs3_4(FloatRegFile_2_io_rs3_4),
    .io_rs3_5(FloatRegFile_2_io_rs3_5),
    .io_rs3_6(FloatRegFile_2_io_rs3_6),
    .io_rs3_7(FloatRegFile_2_io_rs3_7),
    .io_rs1idx(FloatRegFile_2_io_rs1idx),
    .io_rs2idx(FloatRegFile_2_io_rs2idx),
    .io_rs3idx(FloatRegFile_2_io_rs3idx),
    .io_rd_0(FloatRegFile_2_io_rd_0),
    .io_rd_1(FloatRegFile_2_io_rd_1),
    .io_rd_2(FloatRegFile_2_io_rd_2),
    .io_rd_3(FloatRegFile_2_io_rd_3),
    .io_rd_4(FloatRegFile_2_io_rd_4),
    .io_rd_5(FloatRegFile_2_io_rd_5),
    .io_rd_6(FloatRegFile_2_io_rd_6),
    .io_rd_7(FloatRegFile_2_io_rd_7),
    .io_rdidx(FloatRegFile_2_io_rdidx),
    .io_rdwen(FloatRegFile_2_io_rdwen),
    .io_rdwmask_0(FloatRegFile_2_io_rdwmask_0),
    .io_rdwmask_1(FloatRegFile_2_io_rdwmask_1),
    .io_rdwmask_2(FloatRegFile_2_io_rdwmask_2),
    .io_rdwmask_3(FloatRegFile_2_io_rdwmask_3),
    .io_rdwmask_4(FloatRegFile_2_io_rdwmask_4),
    .io_rdwmask_5(FloatRegFile_2_io_rdwmask_5),
    .io_rdwmask_6(FloatRegFile_2_io_rdwmask_6),
    .io_rdwmask_7(FloatRegFile_2_io_rdwmask_7)
  );
  FloatRegFile FloatRegFile_3 ( // @[operandCollector.scala 34:54]
    .clock(FloatRegFile_3_clock),
    .io_v0_0(FloatRegFile_3_io_v0_0),
    .io_rs1_0(FloatRegFile_3_io_rs1_0),
    .io_rs1_1(FloatRegFile_3_io_rs1_1),
    .io_rs1_2(FloatRegFile_3_io_rs1_2),
    .io_rs1_3(FloatRegFile_3_io_rs1_3),
    .io_rs1_4(FloatRegFile_3_io_rs1_4),
    .io_rs1_5(FloatRegFile_3_io_rs1_5),
    .io_rs1_6(FloatRegFile_3_io_rs1_6),
    .io_rs1_7(FloatRegFile_3_io_rs1_7),
    .io_rs2_0(FloatRegFile_3_io_rs2_0),
    .io_rs2_1(FloatRegFile_3_io_rs2_1),
    .io_rs2_2(FloatRegFile_3_io_rs2_2),
    .io_rs2_3(FloatRegFile_3_io_rs2_3),
    .io_rs2_4(FloatRegFile_3_io_rs2_4),
    .io_rs2_5(FloatRegFile_3_io_rs2_5),
    .io_rs2_6(FloatRegFile_3_io_rs2_6),
    .io_rs2_7(FloatRegFile_3_io_rs2_7),
    .io_rs3_0(FloatRegFile_3_io_rs3_0),
    .io_rs3_1(FloatRegFile_3_io_rs3_1),
    .io_rs3_2(FloatRegFile_3_io_rs3_2),
    .io_rs3_3(FloatRegFile_3_io_rs3_3),
    .io_rs3_4(FloatRegFile_3_io_rs3_4),
    .io_rs3_5(FloatRegFile_3_io_rs3_5),
    .io_rs3_6(FloatRegFile_3_io_rs3_6),
    .io_rs3_7(FloatRegFile_3_io_rs3_7),
    .io_rs1idx(FloatRegFile_3_io_rs1idx),
    .io_rs2idx(FloatRegFile_3_io_rs2idx),
    .io_rs3idx(FloatRegFile_3_io_rs3idx),
    .io_rd_0(FloatRegFile_3_io_rd_0),
    .io_rd_1(FloatRegFile_3_io_rd_1),
    .io_rd_2(FloatRegFile_3_io_rd_2),
    .io_rd_3(FloatRegFile_3_io_rd_3),
    .io_rd_4(FloatRegFile_3_io_rd_4),
    .io_rd_5(FloatRegFile_3_io_rd_5),
    .io_rd_6(FloatRegFile_3_io_rd_6),
    .io_rd_7(FloatRegFile_3_io_rd_7),
    .io_rdidx(FloatRegFile_3_io_rdidx),
    .io_rdwen(FloatRegFile_3_io_rdwen),
    .io_rdwmask_0(FloatRegFile_3_io_rdwmask_0),
    .io_rdwmask_1(FloatRegFile_3_io_rdwmask_1),
    .io_rdwmask_2(FloatRegFile_3_io_rdwmask_2),
    .io_rdwmask_3(FloatRegFile_3_io_rdwmask_3),
    .io_rdwmask_4(FloatRegFile_3_io_rdwmask_4),
    .io_rdwmask_5(FloatRegFile_3_io_rdwmask_5),
    .io_rdwmask_6(FloatRegFile_3_io_rdwmask_6),
    .io_rdwmask_7(FloatRegFile_3_io_rdwmask_7)
  );
  RegFile RegFile ( // @[operandCollector.scala 35:54]
    .clock(RegFile_clock),
    .io_rs1(RegFile_io_rs1),
    .io_rs2(RegFile_io_rs2),
    .io_rs3(RegFile_io_rs3),
    .io_rs1idx(RegFile_io_rs1idx),
    .io_rs2idx(RegFile_io_rs2idx),
    .io_rs3idx(RegFile_io_rs3idx),
    .io_rd(RegFile_io_rd),
    .io_rdidx(RegFile_io_rdidx),
    .io_rdwen(RegFile_io_rdwen)
  );
  RegFile RegFile_1 ( // @[operandCollector.scala 35:54]
    .clock(RegFile_1_clock),
    .io_rs1(RegFile_1_io_rs1),
    .io_rs2(RegFile_1_io_rs2),
    .io_rs3(RegFile_1_io_rs3),
    .io_rs1idx(RegFile_1_io_rs1idx),
    .io_rs2idx(RegFile_1_io_rs2idx),
    .io_rs3idx(RegFile_1_io_rs3idx),
    .io_rd(RegFile_1_io_rd),
    .io_rdidx(RegFile_1_io_rdidx),
    .io_rdwen(RegFile_1_io_rdwen)
  );
  RegFile RegFile_2 ( // @[operandCollector.scala 35:54]
    .clock(RegFile_2_clock),
    .io_rs1(RegFile_2_io_rs1),
    .io_rs2(RegFile_2_io_rs2),
    .io_rs3(RegFile_2_io_rs3),
    .io_rs1idx(RegFile_2_io_rs1idx),
    .io_rs2idx(RegFile_2_io_rs2idx),
    .io_rs3idx(RegFile_2_io_rs3idx),
    .io_rd(RegFile_2_io_rd),
    .io_rdidx(RegFile_2_io_rdidx),
    .io_rdwen(RegFile_2_io_rdwen)
  );
  RegFile RegFile_3 ( // @[operandCollector.scala 35:54]
    .clock(RegFile_3_clock),
    .io_rs1(RegFile_3_io_rs1),
    .io_rs2(RegFile_3_io_rs2),
    .io_rs3(RegFile_3_io_rs3),
    .io_rs1idx(RegFile_3_io_rs1idx),
    .io_rs2idx(RegFile_3_io_rs2idx),
    .io_rs3idx(RegFile_3_io_rs3idx),
    .io_rd(RegFile_3_io_rd),
    .io_rdidx(RegFile_3_io_rdidx),
    .io_rdwen(RegFile_3_io_rdwen)
  );
  ImmGen imm ( // @[operandCollector.scala 36:17]
    .io_inst(imm_io_inst),
    .io_sel(imm_io_sel),
    .io_out(imm_io_out)
  );
  assign io_alu_src1_0 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_0_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_1 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_1_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_2 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_2_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_3 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_3_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_4 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_4_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_5 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_5_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_6 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_6_T_3; // @[Mux.scala 81:58]
  assign io_alu_src1_7 = 2'h0 == io_control_sel_alu1 ? io_control_pc : _io_alu_src1_7_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_0 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_0_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_1 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_1_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_2 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_2_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_3 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_3_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_4 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_4_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_5 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_5_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_6 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_6_T_3; // @[Mux.scala 81:58]
  assign io_alu_src2_7 = 2'h0 == io_control_sel_alu2 ? 32'h4 : _io_alu_src2_7_T_3; // @[Mux.scala 81:58]
  assign io_alu_src3_0 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_0_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_1 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_1_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_2 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_2_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_3 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_3_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_4 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_4_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_5 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_5_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_6 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_6_T_10; // @[Mux.scala 81:58]
  assign io_alu_src3_7 = 2'h2 == io_control_sel_alu3 ? _GEN_31 : _io_alu_src3_7_T_10; // @[Mux.scala 81:58]
  assign io_mask_0 = io_control_mask ? _GEN_35[0] : 1'h1; // @[operandCollector.scala 68:20]
  assign io_mask_1 = io_control_mask ? _GEN_35[1] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign io_mask_2 = io_control_mask ? _GEN_35[2] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign io_mask_3 = io_control_mask ? _GEN_35[3] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign io_mask_4 = io_control_mask ? _GEN_35[4] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign io_mask_5 = io_control_mask ? _GEN_35[5] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign io_mask_6 = io_control_mask ? _GEN_35[6] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign io_mask_7 = io_control_mask ? _GEN_35[7] : io_control_isvec; // @[operandCollector.scala 68:20]
  assign FloatRegFile_clock = clock;
  assign FloatRegFile_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 34:28 41:13]
  assign FloatRegFile_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 34:28 42:13]
  assign FloatRegFile_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 34:28 43:13]
  assign FloatRegFile_io_rd_0 = io_writeVecCtrl_bits_wb_wfd_rd_0; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_1 = io_writeVecCtrl_bits_wb_wfd_rd_1; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_2 = io_writeVecCtrl_bits_wb_wfd_rd_2; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_3 = io_writeVecCtrl_bits_wb_wfd_rd_3; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_4 = io_writeVecCtrl_bits_wb_wfd_rd_4; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_5 = io_writeVecCtrl_bits_wb_wfd_rd_5; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_6 = io_writeVecCtrl_bits_wb_wfd_rd_6; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rd_7 = io_writeVecCtrl_bits_wb_wfd_rd_7; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_io_rdidx = io_writeVecCtrl_bits_reg_idxw; // @[operandCollector.scala 34:28 44:12]
  assign FloatRegFile_io_rdwen = 2'h0 == io_writeVecCtrl_bits_warp_id & (io_writeVecCtrl_bits_wfd &
    io_writeVecCtrl_valid); // @[operandCollector.scala 46:12 59:{52,52}]
  assign FloatRegFile_io_rdwmask_0 = io_writeVecCtrl_bits_wfd_mask_0; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_1 = io_writeVecCtrl_bits_wfd_mask_1; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_2 = io_writeVecCtrl_bits_wfd_mask_2; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_3 = io_writeVecCtrl_bits_wfd_mask_3; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_4 = io_writeVecCtrl_bits_wfd_mask_4; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_5 = io_writeVecCtrl_bits_wfd_mask_5; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_6 = io_writeVecCtrl_bits_wfd_mask_6; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_io_rdwmask_7 = io_writeVecCtrl_bits_wfd_mask_7; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_clock = clock;
  assign FloatRegFile_1_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 34:28 41:13]
  assign FloatRegFile_1_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 34:28 42:13]
  assign FloatRegFile_1_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 34:28 43:13]
  assign FloatRegFile_1_io_rd_0 = io_writeVecCtrl_bits_wb_wfd_rd_0; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_1 = io_writeVecCtrl_bits_wb_wfd_rd_1; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_2 = io_writeVecCtrl_bits_wb_wfd_rd_2; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_3 = io_writeVecCtrl_bits_wb_wfd_rd_3; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_4 = io_writeVecCtrl_bits_wb_wfd_rd_4; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_5 = io_writeVecCtrl_bits_wb_wfd_rd_5; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_6 = io_writeVecCtrl_bits_wb_wfd_rd_6; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rd_7 = io_writeVecCtrl_bits_wb_wfd_rd_7; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_1_io_rdidx = io_writeVecCtrl_bits_reg_idxw; // @[operandCollector.scala 34:28 44:12]
  assign FloatRegFile_1_io_rdwen = 2'h1 == io_writeVecCtrl_bits_warp_id & (io_writeVecCtrl_bits_wfd &
    io_writeVecCtrl_valid); // @[operandCollector.scala 46:12 59:{52,52}]
  assign FloatRegFile_1_io_rdwmask_0 = io_writeVecCtrl_bits_wfd_mask_0; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_1 = io_writeVecCtrl_bits_wfd_mask_1; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_2 = io_writeVecCtrl_bits_wfd_mask_2; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_3 = io_writeVecCtrl_bits_wfd_mask_3; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_4 = io_writeVecCtrl_bits_wfd_mask_4; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_5 = io_writeVecCtrl_bits_wfd_mask_5; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_6 = io_writeVecCtrl_bits_wfd_mask_6; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_1_io_rdwmask_7 = io_writeVecCtrl_bits_wfd_mask_7; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_clock = clock;
  assign FloatRegFile_2_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 34:28 41:13]
  assign FloatRegFile_2_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 34:28 42:13]
  assign FloatRegFile_2_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 34:28 43:13]
  assign FloatRegFile_2_io_rd_0 = io_writeVecCtrl_bits_wb_wfd_rd_0; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_1 = io_writeVecCtrl_bits_wb_wfd_rd_1; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_2 = io_writeVecCtrl_bits_wb_wfd_rd_2; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_3 = io_writeVecCtrl_bits_wb_wfd_rd_3; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_4 = io_writeVecCtrl_bits_wb_wfd_rd_4; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_5 = io_writeVecCtrl_bits_wb_wfd_rd_5; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_6 = io_writeVecCtrl_bits_wb_wfd_rd_6; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rd_7 = io_writeVecCtrl_bits_wb_wfd_rd_7; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_2_io_rdidx = io_writeVecCtrl_bits_reg_idxw; // @[operandCollector.scala 34:28 44:12]
  assign FloatRegFile_2_io_rdwen = 2'h2 == io_writeVecCtrl_bits_warp_id & (io_writeVecCtrl_bits_wfd &
    io_writeVecCtrl_valid); // @[operandCollector.scala 46:12 59:{52,52}]
  assign FloatRegFile_2_io_rdwmask_0 = io_writeVecCtrl_bits_wfd_mask_0; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_1 = io_writeVecCtrl_bits_wfd_mask_1; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_2 = io_writeVecCtrl_bits_wfd_mask_2; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_3 = io_writeVecCtrl_bits_wfd_mask_3; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_4 = io_writeVecCtrl_bits_wfd_mask_4; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_5 = io_writeVecCtrl_bits_wfd_mask_5; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_6 = io_writeVecCtrl_bits_wfd_mask_6; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_2_io_rdwmask_7 = io_writeVecCtrl_bits_wfd_mask_7; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_clock = clock;
  assign FloatRegFile_3_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 34:28 41:13]
  assign FloatRegFile_3_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 34:28 42:13]
  assign FloatRegFile_3_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 34:28 43:13]
  assign FloatRegFile_3_io_rd_0 = io_writeVecCtrl_bits_wb_wfd_rd_0; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_1 = io_writeVecCtrl_bits_wb_wfd_rd_1; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_2 = io_writeVecCtrl_bits_wb_wfd_rd_2; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_3 = io_writeVecCtrl_bits_wb_wfd_rd_3; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_4 = io_writeVecCtrl_bits_wb_wfd_rd_4; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_5 = io_writeVecCtrl_bits_wb_wfd_rd_5; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_6 = io_writeVecCtrl_bits_wb_wfd_rd_6; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rd_7 = io_writeVecCtrl_bits_wb_wfd_rd_7; // @[operandCollector.scala 34:28 45:9]
  assign FloatRegFile_3_io_rdidx = io_writeVecCtrl_bits_reg_idxw; // @[operandCollector.scala 34:28 44:12]
  assign FloatRegFile_3_io_rdwen = 2'h3 == io_writeVecCtrl_bits_warp_id & (io_writeVecCtrl_bits_wfd &
    io_writeVecCtrl_valid); // @[operandCollector.scala 46:12 59:{52,52}]
  assign FloatRegFile_3_io_rdwmask_0 = io_writeVecCtrl_bits_wfd_mask_0; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_1 = io_writeVecCtrl_bits_wfd_mask_1; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_2 = io_writeVecCtrl_bits_wfd_mask_2; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_3 = io_writeVecCtrl_bits_wfd_mask_3; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_4 = io_writeVecCtrl_bits_wfd_mask_4; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_5 = io_writeVecCtrl_bits_wfd_mask_5; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_6 = io_writeVecCtrl_bits_wfd_mask_6; // @[operandCollector.scala 34:28 47:14]
  assign FloatRegFile_3_io_rdwmask_7 = io_writeVecCtrl_bits_wfd_mask_7; // @[operandCollector.scala 34:28 47:14]
  assign RegFile_clock = clock;
  assign RegFile_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 35:28 51:13]
  assign RegFile_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 35:28 52:13]
  assign RegFile_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 35:28 53:13]
  assign RegFile_io_rd = io_writeScalarCtrl_bits_wb_wxd_rd; // @[operandCollector.scala 35:28 55:9]
  assign RegFile_io_rdidx = io_writeScalarCtrl_bits_reg_idxw; // @[operandCollector.scala 35:28 54:12]
  assign RegFile_io_rdwen = 2'h0 == io_writeScalarCtrl_bits_warp_id & (io_writeScalarCtrl_bits_wxd &
    io_writeScalarCtrl_valid); // @[operandCollector.scala 56:12 60:{55,55}]
  assign RegFile_1_clock = clock;
  assign RegFile_1_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 35:28 51:13]
  assign RegFile_1_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 35:28 52:13]
  assign RegFile_1_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 35:28 53:13]
  assign RegFile_1_io_rd = io_writeScalarCtrl_bits_wb_wxd_rd; // @[operandCollector.scala 35:28 55:9]
  assign RegFile_1_io_rdidx = io_writeScalarCtrl_bits_reg_idxw; // @[operandCollector.scala 35:28 54:12]
  assign RegFile_1_io_rdwen = 2'h1 == io_writeScalarCtrl_bits_warp_id & (io_writeScalarCtrl_bits_wxd &
    io_writeScalarCtrl_valid); // @[operandCollector.scala 56:12 60:{55,55}]
  assign RegFile_2_clock = clock;
  assign RegFile_2_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 35:28 51:13]
  assign RegFile_2_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 35:28 52:13]
  assign RegFile_2_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 35:28 53:13]
  assign RegFile_2_io_rd = io_writeScalarCtrl_bits_wb_wxd_rd; // @[operandCollector.scala 35:28 55:9]
  assign RegFile_2_io_rdidx = io_writeScalarCtrl_bits_reg_idxw; // @[operandCollector.scala 35:28 54:12]
  assign RegFile_2_io_rdwen = 2'h2 == io_writeScalarCtrl_bits_warp_id & (io_writeScalarCtrl_bits_wxd &
    io_writeScalarCtrl_valid); // @[operandCollector.scala 56:12 60:{55,55}]
  assign RegFile_3_clock = clock;
  assign RegFile_3_io_rs1idx = io_control_reg_idx1; // @[operandCollector.scala 35:28 51:13]
  assign RegFile_3_io_rs2idx = io_control_reg_idx2; // @[operandCollector.scala 35:28 52:13]
  assign RegFile_3_io_rs3idx = io_control_reg_idx3; // @[operandCollector.scala 35:28 53:13]
  assign RegFile_3_io_rd = io_writeScalarCtrl_bits_wb_wxd_rd; // @[operandCollector.scala 35:28 55:9]
  assign RegFile_3_io_rdidx = io_writeScalarCtrl_bits_reg_idxw; // @[operandCollector.scala 35:28 54:12]
  assign RegFile_3_io_rdwen = 2'h3 == io_writeScalarCtrl_bits_warp_id & (io_writeScalarCtrl_bits_wxd &
    io_writeScalarCtrl_valid); // @[operandCollector.scala 56:12 60:{55,55}]
  assign imm_io_inst = io_control_inst; // @[operandCollector.scala 37:14]
  assign imm_io_sel = io_control_sel_imm; // @[operandCollector.scala 38:13]
endmodule
module Issue(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_in1_0,
  input  [31:0] io_in_bits_in1_1,
  input  [31:0] io_in_bits_in1_2,
  input  [31:0] io_in_bits_in1_3,
  input  [31:0] io_in_bits_in1_4,
  input  [31:0] io_in_bits_in1_5,
  input  [31:0] io_in_bits_in1_6,
  input  [31:0] io_in_bits_in1_7,
  input  [31:0] io_in_bits_in2_0,
  input  [31:0] io_in_bits_in2_1,
  input  [31:0] io_in_bits_in2_2,
  input  [31:0] io_in_bits_in2_3,
  input  [31:0] io_in_bits_in2_4,
  input  [31:0] io_in_bits_in2_5,
  input  [31:0] io_in_bits_in2_6,
  input  [31:0] io_in_bits_in2_7,
  input  [31:0] io_in_bits_in3_0,
  input  [31:0] io_in_bits_in3_1,
  input  [31:0] io_in_bits_in3_2,
  input  [31:0] io_in_bits_in3_3,
  input  [31:0] io_in_bits_in3_4,
  input  [31:0] io_in_bits_in3_5,
  input  [31:0] io_in_bits_in3_6,
  input  [31:0] io_in_bits_in3_7,
  input         io_in_bits_mask_0,
  input         io_in_bits_mask_1,
  input         io_in_bits_mask_2,
  input         io_in_bits_mask_3,
  input         io_in_bits_mask_4,
  input         io_in_bits_mask_5,
  input         io_in_bits_mask_6,
  input         io_in_bits_mask_7,
  input  [31:0] io_in_bits_ctrl_inst,
  input  [1:0]  io_in_bits_ctrl_wid,
  input         io_in_bits_ctrl_fp,
  input  [1:0]  io_in_bits_ctrl_branch,
  input         io_in_bits_ctrl_simt_stack,
  input         io_in_bits_ctrl_simt_stack_op,
  input         io_in_bits_ctrl_barrier,
  input  [1:0]  io_in_bits_ctrl_csr,
  input         io_in_bits_ctrl_reverse,
  input         io_in_bits_ctrl_isvec,
  input         io_in_bits_ctrl_mem_unsigned,
  input  [5:0]  io_in_bits_ctrl_alu_fn,
  input         io_in_bits_ctrl_mem,
  input  [1:0]  io_in_bits_ctrl_mem_cmd,
  input  [1:0]  io_in_bits_ctrl_mop,
  input  [4:0]  io_in_bits_ctrl_reg_idxw,
  input         io_in_bits_ctrl_wfd,
  input         io_in_bits_ctrl_fence,
  input         io_in_bits_ctrl_sfu,
  input         io_in_bits_ctrl_readmask,
  input         io_in_bits_ctrl_writemask,
  input         io_in_bits_ctrl_wxd,
  input  [31:0] io_in_bits_ctrl_pc,
  input         io_out_sALU_ready,
  output        io_out_sALU_valid,
  output [31:0] io_out_sALU_bits_in1,
  output [31:0] io_out_sALU_bits_in2,
  output [31:0] io_out_sALU_bits_in3,
  output [1:0]  io_out_sALU_bits_ctrl_wid,
  output [1:0]  io_out_sALU_bits_ctrl_branch,
  output [5:0]  io_out_sALU_bits_ctrl_alu_fn,
  output [4:0]  io_out_sALU_bits_ctrl_reg_idxw,
  output        io_out_sALU_bits_ctrl_wxd,
  input         io_out_vALU_ready,
  output        io_out_vALU_valid,
  output [31:0] io_out_vALU_bits_in1_0,
  output [31:0] io_out_vALU_bits_in1_1,
  output [31:0] io_out_vALU_bits_in1_2,
  output [31:0] io_out_vALU_bits_in1_3,
  output [31:0] io_out_vALU_bits_in1_4,
  output [31:0] io_out_vALU_bits_in1_5,
  output [31:0] io_out_vALU_bits_in1_6,
  output [31:0] io_out_vALU_bits_in1_7,
  output [31:0] io_out_vALU_bits_in2_0,
  output [31:0] io_out_vALU_bits_in2_1,
  output [31:0] io_out_vALU_bits_in2_2,
  output [31:0] io_out_vALU_bits_in2_3,
  output [31:0] io_out_vALU_bits_in2_4,
  output [31:0] io_out_vALU_bits_in2_5,
  output [31:0] io_out_vALU_bits_in2_6,
  output [31:0] io_out_vALU_bits_in2_7,
  output [31:0] io_out_vALU_bits_in3_0,
  output [31:0] io_out_vALU_bits_in3_1,
  output [31:0] io_out_vALU_bits_in3_2,
  output [31:0] io_out_vALU_bits_in3_3,
  output [31:0] io_out_vALU_bits_in3_4,
  output [31:0] io_out_vALU_bits_in3_5,
  output [31:0] io_out_vALU_bits_in3_6,
  output [31:0] io_out_vALU_bits_in3_7,
  output        io_out_vALU_bits_mask_0,
  output        io_out_vALU_bits_mask_1,
  output        io_out_vALU_bits_mask_2,
  output        io_out_vALU_bits_mask_3,
  output        io_out_vALU_bits_mask_4,
  output        io_out_vALU_bits_mask_5,
  output        io_out_vALU_bits_mask_6,
  output        io_out_vALU_bits_mask_7,
  output [1:0]  io_out_vALU_bits_ctrl_wid,
  output        io_out_vALU_bits_ctrl_simt_stack,
  output        io_out_vALU_bits_ctrl_reverse,
  output [5:0]  io_out_vALU_bits_ctrl_alu_fn,
  output [4:0]  io_out_vALU_bits_ctrl_reg_idxw,
  output        io_out_vALU_bits_ctrl_wfd,
  output        io_out_vALU_bits_ctrl_readmask,
  output        io_out_vALU_bits_ctrl_writemask,
  input         io_out_vFPU_ready,
  output        io_out_vFPU_valid,
  output [31:0] io_out_vFPU_bits_in1_0,
  output [31:0] io_out_vFPU_bits_in1_1,
  output [31:0] io_out_vFPU_bits_in1_2,
  output [31:0] io_out_vFPU_bits_in1_3,
  output [31:0] io_out_vFPU_bits_in1_4,
  output [31:0] io_out_vFPU_bits_in1_5,
  output [31:0] io_out_vFPU_bits_in1_6,
  output [31:0] io_out_vFPU_bits_in1_7,
  output [31:0] io_out_vFPU_bits_in2_0,
  output [31:0] io_out_vFPU_bits_in2_1,
  output [31:0] io_out_vFPU_bits_in2_2,
  output [31:0] io_out_vFPU_bits_in2_3,
  output [31:0] io_out_vFPU_bits_in2_4,
  output [31:0] io_out_vFPU_bits_in2_5,
  output [31:0] io_out_vFPU_bits_in2_6,
  output [31:0] io_out_vFPU_bits_in2_7,
  output [31:0] io_out_vFPU_bits_in3_0,
  output [31:0] io_out_vFPU_bits_in3_1,
  output [31:0] io_out_vFPU_bits_in3_2,
  output [31:0] io_out_vFPU_bits_in3_3,
  output [31:0] io_out_vFPU_bits_in3_4,
  output [31:0] io_out_vFPU_bits_in3_5,
  output [31:0] io_out_vFPU_bits_in3_6,
  output [31:0] io_out_vFPU_bits_in3_7,
  output        io_out_vFPU_bits_mask_0,
  output        io_out_vFPU_bits_mask_1,
  output        io_out_vFPU_bits_mask_2,
  output        io_out_vFPU_bits_mask_3,
  output        io_out_vFPU_bits_mask_4,
  output        io_out_vFPU_bits_mask_5,
  output        io_out_vFPU_bits_mask_6,
  output        io_out_vFPU_bits_mask_7,
  output [1:0]  io_out_vFPU_bits_ctrl_wid,
  output        io_out_vFPU_bits_ctrl_reverse,
  output [5:0]  io_out_vFPU_bits_ctrl_alu_fn,
  output [4:0]  io_out_vFPU_bits_ctrl_reg_idxw,
  output        io_out_vFPU_bits_ctrl_wfd,
  output        io_out_vFPU_bits_ctrl_wxd,
  input         io_out_LSU_ready,
  output        io_out_LSU_valid,
  output [31:0] io_out_LSU_bits_in1_0,
  output [31:0] io_out_LSU_bits_in1_1,
  output [31:0] io_out_LSU_bits_in1_2,
  output [31:0] io_out_LSU_bits_in1_3,
  output [31:0] io_out_LSU_bits_in1_4,
  output [31:0] io_out_LSU_bits_in1_5,
  output [31:0] io_out_LSU_bits_in1_6,
  output [31:0] io_out_LSU_bits_in1_7,
  output [31:0] io_out_LSU_bits_in2_0,
  output [31:0] io_out_LSU_bits_in2_1,
  output [31:0] io_out_LSU_bits_in2_2,
  output [31:0] io_out_LSU_bits_in2_3,
  output [31:0] io_out_LSU_bits_in2_4,
  output [31:0] io_out_LSU_bits_in2_5,
  output [31:0] io_out_LSU_bits_in2_6,
  output [31:0] io_out_LSU_bits_in2_7,
  output [31:0] io_out_LSU_bits_in3_0,
  output [31:0] io_out_LSU_bits_in3_1,
  output [31:0] io_out_LSU_bits_in3_2,
  output [31:0] io_out_LSU_bits_in3_3,
  output [31:0] io_out_LSU_bits_in3_4,
  output [31:0] io_out_LSU_bits_in3_5,
  output [31:0] io_out_LSU_bits_in3_6,
  output [31:0] io_out_LSU_bits_in3_7,
  output        io_out_LSU_bits_mask_0,
  output        io_out_LSU_bits_mask_1,
  output        io_out_LSU_bits_mask_2,
  output        io_out_LSU_bits_mask_3,
  output        io_out_LSU_bits_mask_4,
  output        io_out_LSU_bits_mask_5,
  output        io_out_LSU_bits_mask_6,
  output        io_out_LSU_bits_mask_7,
  output [31:0] io_out_LSU_bits_ctrl_inst,
  output [1:0]  io_out_LSU_bits_ctrl_wid,
  output        io_out_LSU_bits_ctrl_fp,
  output [1:0]  io_out_LSU_bits_ctrl_branch,
  output        io_out_LSU_bits_ctrl_simt_stack,
  output        io_out_LSU_bits_ctrl_simt_stack_op,
  output        io_out_LSU_bits_ctrl_barrier,
  output [1:0]  io_out_LSU_bits_ctrl_csr,
  output        io_out_LSU_bits_ctrl_reverse,
  output        io_out_LSU_bits_ctrl_isvec,
  output        io_out_LSU_bits_ctrl_mem_unsigned,
  output [5:0]  io_out_LSU_bits_ctrl_alu_fn,
  output        io_out_LSU_bits_ctrl_mem,
  output [1:0]  io_out_LSU_bits_ctrl_mem_cmd,
  output [1:0]  io_out_LSU_bits_ctrl_mop,
  output [4:0]  io_out_LSU_bits_ctrl_reg_idxw,
  output        io_out_LSU_bits_ctrl_wfd,
  output        io_out_LSU_bits_ctrl_fence,
  output        io_out_LSU_bits_ctrl_sfu,
  output        io_out_LSU_bits_ctrl_readmask,
  output        io_out_LSU_bits_ctrl_writemask,
  output        io_out_LSU_bits_ctrl_wxd,
  output [31:0] io_out_LSU_bits_ctrl_pc,
  input         io_out_SFU_ready,
  output        io_out_SFU_valid,
  output [31:0] io_out_SFU_bits_in1_0,
  output [31:0] io_out_SFU_bits_in1_1,
  output [31:0] io_out_SFU_bits_in1_2,
  output [31:0] io_out_SFU_bits_in1_3,
  output [31:0] io_out_SFU_bits_in1_4,
  output [31:0] io_out_SFU_bits_in1_5,
  output [31:0] io_out_SFU_bits_in1_6,
  output [31:0] io_out_SFU_bits_in1_7,
  output [31:0] io_out_SFU_bits_in2_0,
  output [31:0] io_out_SFU_bits_in2_1,
  output [31:0] io_out_SFU_bits_in2_2,
  output [31:0] io_out_SFU_bits_in2_3,
  output [31:0] io_out_SFU_bits_in2_4,
  output [31:0] io_out_SFU_bits_in2_5,
  output [31:0] io_out_SFU_bits_in2_6,
  output [31:0] io_out_SFU_bits_in2_7,
  output        io_out_SFU_bits_mask_0,
  output        io_out_SFU_bits_mask_1,
  output        io_out_SFU_bits_mask_2,
  output        io_out_SFU_bits_mask_3,
  output        io_out_SFU_bits_mask_4,
  output        io_out_SFU_bits_mask_5,
  output        io_out_SFU_bits_mask_6,
  output        io_out_SFU_bits_mask_7,
  output [1:0]  io_out_SFU_bits_ctrl_wid,
  output        io_out_SFU_bits_ctrl_fp,
  output        io_out_SFU_bits_ctrl_reverse,
  output        io_out_SFU_bits_ctrl_isvec,
  output [5:0]  io_out_SFU_bits_ctrl_alu_fn,
  output [4:0]  io_out_SFU_bits_ctrl_reg_idxw,
  output        io_out_SFU_bits_ctrl_wfd,
  output        io_out_SFU_bits_ctrl_wxd,
  input         io_out_SIMT_ready,
  output        io_out_SIMT_valid,
  output        io_out_SIMT_bits_opcode,
  output [1:0]  io_out_SIMT_bits_wid,
  output [31:0] io_out_SIMT_bits_PC_branch,
  output [7:0]  io_out_SIMT_bits_mask_init,
  input         io_out_warpscheduler_ready,
  output        io_out_warpscheduler_valid,
  output [1:0]  io_out_warpscheduler_bits_ctrl_wid,
  output        io_out_warpscheduler_bits_ctrl_simt_stack_op,
  output        io_out_warpscheduler_bits_ctrl_barrier,
  input         io_out_CSR_ready,
  output        io_out_CSR_valid,
  output [31:0] io_out_CSR_bits_ctrl_inst,
  output [1:0]  io_out_CSR_bits_ctrl_wid,
  output [1:0]  io_out_CSR_bits_ctrl_csr,
  output        io_out_CSR_bits_ctrl_isvec,
  output [4:0]  io_out_CSR_bits_ctrl_reg_idxw,
  output        io_out_CSR_bits_ctrl_wxd,
  output [31:0] io_out_CSR_bits_in1
);
  wire [3:0] io_out_SIMT_bits_mask_init_lo = {io_in_bits_mask_3,io_in_bits_mask_2,io_in_bits_mask_1,io_in_bits_mask_0}; // @[issue.scala 56:56]
  wire [3:0] io_out_SIMT_bits_mask_init_hi = {io_in_bits_mask_7,io_in_bits_mask_6,io_in_bits_mask_5,io_in_bits_mask_4}; // @[issue.scala 56:56]
  wire  beqv_ready = io_out_SIMT_ready & io_out_vALU_ready; // @[issue.scala 88:39]
  wire  _io_out_vALU_valid_T = io_in_valid & beqv_ready; // @[issue.scala 89:41]
  wire  _GEN_0 = ~io_out_SIMT_bits_opcode & (io_in_valid & beqv_ready); // @[issue.scala 63:20 87:44 89:24]
  wire  _GEN_1 = ~io_out_SIMT_bits_opcode ? _io_out_vALU_valid_T : io_in_valid; // @[issue.scala 87:44 90:24 93:26]
  wire  _GEN_2 = ~io_out_SIMT_bits_opcode ? beqv_ready : io_out_SIMT_ready; // @[issue.scala 87:44 91:21 94:23]
  wire  _GEN_3 = io_in_bits_ctrl_simt_stack ? _GEN_0 : io_in_valid; // @[issue.scala 86:40 97:24]
  wire  _GEN_4 = io_in_bits_ctrl_simt_stack & _GEN_1; // @[issue.scala 64:20 86:40]
  wire  _GEN_5 = io_in_bits_ctrl_simt_stack ? _GEN_2 : io_out_vALU_ready; // @[issue.scala 86:40 98:21]
  wire  _GEN_6 = io_in_bits_ctrl_barrier & io_in_valid; // @[issue.scala 100:41 101:31 67:29]
  wire  _GEN_7 = io_in_bits_ctrl_barrier ? io_out_warpscheduler_ready : io_out_sALU_ready; // @[issue.scala 100:41 102:19 105:19]
  wire  _GEN_8 = io_in_bits_ctrl_barrier ? 1'h0 : io_in_valid; // @[issue.scala 100:41 62:20 104:22]
  wire  _GEN_9 = io_in_bits_ctrl_isvec & _GEN_3; // @[issue.scala 63:20 85:39]
  wire  _GEN_10 = io_in_bits_ctrl_isvec & _GEN_4; // @[issue.scala 64:20 85:39]
  wire  _GEN_11 = io_in_bits_ctrl_isvec ? _GEN_5 : _GEN_7; // @[issue.scala 85:39]
  wire  _GEN_12 = io_in_bits_ctrl_isvec ? 1'h0 : _GEN_6; // @[issue.scala 67:29 85:39]
  wire  _GEN_13 = io_in_bits_ctrl_isvec ? 1'h0 : _GEN_8; // @[issue.scala 62:20 85:39]
  wire  _GEN_14 = io_in_bits_ctrl_mem & io_in_valid; // @[issue.scala 65:19 81:38 83:21]
  wire  _GEN_15 = io_in_bits_ctrl_mem ? io_out_LSU_ready : _GEN_11; // @[issue.scala 81:38 84:19]
  wire  _GEN_16 = io_in_bits_ctrl_mem ? 1'h0 : _GEN_9; // @[issue.scala 63:20 81:38]
  wire  _GEN_17 = io_in_bits_ctrl_mem ? 1'h0 : _GEN_10; // @[issue.scala 64:20 81:38]
  wire  _GEN_18 = io_in_bits_ctrl_mem ? 1'h0 : _GEN_12; // @[issue.scala 67:29 81:38]
  wire  _GEN_19 = io_in_bits_ctrl_mem ? 1'h0 : _GEN_13; // @[issue.scala 62:20 81:38]
  wire  _GEN_20 = |io_in_bits_ctrl_csr & io_in_valid; // @[issue.scala 68:19 77:43 78:21]
  wire  _GEN_21 = |io_in_bits_ctrl_csr ? io_out_CSR_ready : _GEN_15; // @[issue.scala 77:43 79:19]
  wire  _GEN_22 = |io_in_bits_ctrl_csr ? 1'h0 : _GEN_14; // @[issue.scala 65:19 77:43]
  wire  _GEN_23 = |io_in_bits_ctrl_csr ? 1'h0 : _GEN_16; // @[issue.scala 63:20 77:43]
  wire  _GEN_24 = |io_in_bits_ctrl_csr ? 1'h0 : _GEN_17; // @[issue.scala 64:20 77:43]
  wire  _GEN_25 = |io_in_bits_ctrl_csr ? 1'h0 : _GEN_18; // @[issue.scala 67:29 77:43]
  wire  _GEN_26 = |io_in_bits_ctrl_csr ? 1'h0 : _GEN_19; // @[issue.scala 62:20 77:43]
  wire  _GEN_27 = io_in_bits_ctrl_fp & io_in_valid; // @[issue.scala 66:20 74:36 75:22]
  wire  _GEN_28 = io_in_bits_ctrl_fp ? io_out_vFPU_ready : _GEN_21; // @[issue.scala 74:36 76:19]
  wire  _GEN_29 = io_in_bits_ctrl_fp ? 1'h0 : _GEN_20; // @[issue.scala 68:19 74:36]
  wire  _GEN_30 = io_in_bits_ctrl_fp ? 1'h0 : _GEN_22; // @[issue.scala 65:19 74:36]
  wire  _GEN_31 = io_in_bits_ctrl_fp ? 1'h0 : _GEN_23; // @[issue.scala 63:20 74:36]
  wire  _GEN_32 = io_in_bits_ctrl_fp ? 1'h0 : _GEN_24; // @[issue.scala 64:20 74:36]
  wire  _GEN_33 = io_in_bits_ctrl_fp ? 1'h0 : _GEN_25; // @[issue.scala 67:29 74:36]
  wire  _GEN_34 = io_in_bits_ctrl_fp ? 1'h0 : _GEN_26; // @[issue.scala 62:20 74:36]
  assign io_in_ready = io_in_bits_ctrl_sfu ? io_out_SFU_ready : _GEN_28; // @[issue.scala 71:31 73:19]
  assign io_out_sALU_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_34; // @[issue.scala 62:20 71:31]
  assign io_out_sALU_bits_in1 = io_in_bits_in1_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_in2 = io_in_bits_in2_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_in3 = io_in_bits_in3_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_ctrl_branch = io_in_bits_ctrl_branch; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_ctrl_alu_fn = io_in_bits_ctrl_alu_fn; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign io_out_sALU_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_31; // @[issue.scala 63:20 71:31]
  assign io_out_vALU_bits_in1_0 = io_in_bits_in1_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_1 = io_in_bits_in1_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_2 = io_in_bits_in1_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_3 = io_in_bits_in1_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_4 = io_in_bits_in1_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_5 = io_in_bits_in1_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_6 = io_in_bits_in1_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in1_7 = io_in_bits_in1_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_0 = io_in_bits_in2_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_1 = io_in_bits_in2_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_2 = io_in_bits_in2_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_3 = io_in_bits_in2_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_4 = io_in_bits_in2_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_5 = io_in_bits_in2_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_6 = io_in_bits_in2_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in2_7 = io_in_bits_in2_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_0 = io_in_bits_in3_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_1 = io_in_bits_in3_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_2 = io_in_bits_in3_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_3 = io_in_bits_in3_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_4 = io_in_bits_in3_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_5 = io_in_bits_in3_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_6 = io_in_bits_in3_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_in3_7 = io_in_bits_in3_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_0 = io_in_bits_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_1 = io_in_bits_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_2 = io_in_bits_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_3 = io_in_bits_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_4 = io_in_bits_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_5 = io_in_bits_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_6 = io_in_bits_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_mask_7 = io_in_bits_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_simt_stack = io_in_bits_ctrl_simt_stack; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_reverse = io_in_bits_ctrl_reverse; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_alu_fn = io_in_bits_ctrl_alu_fn; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_readmask = io_in_bits_ctrl_readmask; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vALU_bits_ctrl_writemask = io_in_bits_ctrl_writemask; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_27; // @[issue.scala 66:20 71:31]
  assign io_out_vFPU_bits_in1_0 = io_in_bits_in1_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_1 = io_in_bits_in1_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_2 = io_in_bits_in1_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_3 = io_in_bits_in1_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_4 = io_in_bits_in1_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_5 = io_in_bits_in1_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_6 = io_in_bits_in1_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in1_7 = io_in_bits_in1_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_0 = io_in_bits_in2_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_1 = io_in_bits_in2_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_2 = io_in_bits_in2_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_3 = io_in_bits_in2_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_4 = io_in_bits_in2_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_5 = io_in_bits_in2_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_6 = io_in_bits_in2_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in2_7 = io_in_bits_in2_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_0 = io_in_bits_in3_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_1 = io_in_bits_in3_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_2 = io_in_bits_in3_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_3 = io_in_bits_in3_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_4 = io_in_bits_in3_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_5 = io_in_bits_in3_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_6 = io_in_bits_in3_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_in3_7 = io_in_bits_in3_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_0 = io_in_bits_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_1 = io_in_bits_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_2 = io_in_bits_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_3 = io_in_bits_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_4 = io_in_bits_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_5 = io_in_bits_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_6 = io_in_bits_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_mask_7 = io_in_bits_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_ctrl_reverse = io_in_bits_ctrl_reverse; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_ctrl_alu_fn = io_in_bits_ctrl_alu_fn; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_vFPU_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_30; // @[issue.scala 65:19 71:31]
  assign io_out_LSU_bits_in1_0 = io_in_bits_in1_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_1 = io_in_bits_in1_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_2 = io_in_bits_in1_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_3 = io_in_bits_in1_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_4 = io_in_bits_in1_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_5 = io_in_bits_in1_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_6 = io_in_bits_in1_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in1_7 = io_in_bits_in1_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_0 = io_in_bits_in2_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_1 = io_in_bits_in2_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_2 = io_in_bits_in2_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_3 = io_in_bits_in2_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_4 = io_in_bits_in2_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_5 = io_in_bits_in2_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_6 = io_in_bits_in2_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in2_7 = io_in_bits_in2_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_0 = io_in_bits_in3_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_1 = io_in_bits_in3_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_2 = io_in_bits_in3_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_3 = io_in_bits_in3_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_4 = io_in_bits_in3_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_5 = io_in_bits_in3_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_6 = io_in_bits_in3_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_in3_7 = io_in_bits_in3_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_0 = io_in_bits_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_1 = io_in_bits_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_2 = io_in_bits_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_3 = io_in_bits_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_4 = io_in_bits_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_5 = io_in_bits_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_6 = io_in_bits_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_mask_7 = io_in_bits_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_inst = io_in_bits_ctrl_inst; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_fp = io_in_bits_ctrl_fp; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_branch = io_in_bits_ctrl_branch; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_simt_stack = io_in_bits_ctrl_simt_stack; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_simt_stack_op = io_in_bits_ctrl_simt_stack_op; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_barrier = io_in_bits_ctrl_barrier; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_csr = io_in_bits_ctrl_csr; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_reverse = io_in_bits_ctrl_reverse; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_isvec = io_in_bits_ctrl_isvec; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_mem_unsigned = io_in_bits_ctrl_mem_unsigned; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_alu_fn = io_in_bits_ctrl_alu_fn; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_mem = io_in_bits_ctrl_mem; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_mem_cmd = io_in_bits_ctrl_mem_cmd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_mop = io_in_bits_ctrl_mop; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_fence = io_in_bits_ctrl_fence; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_sfu = io_in_bits_ctrl_sfu; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_readmask = io_in_bits_ctrl_readmask; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_writemask = io_in_bits_ctrl_writemask; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_LSU_bits_ctrl_pc = io_in_bits_ctrl_pc; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_valid = io_in_bits_ctrl_sfu & io_in_valid; // @[issue.scala 69:19 71:31 72:21]
  assign io_out_SFU_bits_in1_0 = io_in_bits_in1_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_1 = io_in_bits_in1_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_2 = io_in_bits_in1_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_3 = io_in_bits_in1_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_4 = io_in_bits_in1_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_5 = io_in_bits_in1_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_6 = io_in_bits_in1_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in1_7 = io_in_bits_in1_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_0 = io_in_bits_in2_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_1 = io_in_bits_in2_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_2 = io_in_bits_in2_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_3 = io_in_bits_in2_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_4 = io_in_bits_in2_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_5 = io_in_bits_in2_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_6 = io_in_bits_in2_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_in2_7 = io_in_bits_in2_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_0 = io_in_bits_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_1 = io_in_bits_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_2 = io_in_bits_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_3 = io_in_bits_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_4 = io_in_bits_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_5 = io_in_bits_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_6 = io_in_bits_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_mask_7 = io_in_bits_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_fp = io_in_bits_ctrl_fp; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_reverse = io_in_bits_ctrl_reverse; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_isvec = io_in_bits_ctrl_isvec; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_alu_fn = io_in_bits_ctrl_alu_fn; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SFU_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SIMT_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_32; // @[issue.scala 64:20 71:31]
  assign io_out_SIMT_bits_opcode = io_in_bits_ctrl_simt_stack_op; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SIMT_bits_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SIMT_bits_PC_branch = io_in_bits_in3_0; // @[Decoupled.scala 355:21 357:16]
  assign io_out_SIMT_bits_mask_init = {io_out_SIMT_bits_mask_init_hi,io_out_SIMT_bits_mask_init_lo}; // @[issue.scala 56:56]
  assign io_out_warpscheduler_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_33; // @[issue.scala 67:29 71:31]
  assign io_out_warpscheduler_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_warpscheduler_bits_ctrl_simt_stack_op = io_in_bits_ctrl_simt_stack_op; // @[Decoupled.scala 355:21 357:16]
  assign io_out_warpscheduler_bits_ctrl_barrier = io_in_bits_ctrl_barrier; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_valid = io_in_bits_ctrl_sfu ? 1'h0 : _GEN_29; // @[issue.scala 68:19 71:31]
  assign io_out_CSR_bits_ctrl_inst = io_in_bits_ctrl_inst; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_bits_ctrl_csr = io_in_bits_ctrl_csr; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_bits_ctrl_isvec = io_in_bits_ctrl_isvec; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[Decoupled.scala 355:21 357:16]
  assign io_out_CSR_bits_in1 = io_in_bits_in1_0; // @[Decoupled.scala 355:21 357:16]
endmodule
module ScalarALU(
  input  [4:0]  io_func,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  input  [31:0] io_in3,
  output [31:0] io_out,
  output        io_cmp_out
);
  wire  _in2_inv_T_1 = io_func <= 5'hf; // @[ALU.scala 45:49]
  wire  _in2_inv_T_2 = io_func >= 5'ha & io_func <= 5'hf; // @[ALU.scala 45:42]
  wire [31:0] _in2_inv_T_3 = ~io_in2; // @[ALU.scala 69:38]
  wire [31:0] in2_inv = _in2_inv_T_2 ? _in2_inv_T_3 : io_in2; // @[ALU.scala 69:20]
  wire [31:0] _adder_out_T_1 = io_in1 + in2_inv; // @[ALU.scala 70:26]
  wire [31:0] _GEN_0 = {{31'd0}, _in2_inv_T_2}; // @[ALU.scala 70:36]
  wire [31:0] adder_out = _adder_out_T_1 + _GEN_0; // @[ALU.scala 70:36]
  wire [31:0] in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 71:28]
  wire  _slt_T_7 = io_func[1] ? io_in2[31] : io_in1[31]; // @[ALU.scala 76:10]
  wire  slt = io_in1[31] == io_in2[31] ? adder_out[31] : _slt_T_7; // @[ALU.scala 75:8]
  wire  _io_cmp_out_T_2 = ~io_func[3]; // @[ALU.scala 49:26]
  wire  _io_cmp_out_T_4 = _io_cmp_out_T_2 ? in1_xor_in2 == 32'h0 : slt; // @[ALU.scala 77:43]
  wire [4:0] shamt = io_in2[4:0]; // @[ALU.scala 80:32]
  wire  _shin_T_2 = io_func == 5'h5 | io_func == 5'hb; // @[ALU.scala 81:36]
  wire [31:0] _GEN_1 = {{16'd0}, io_in1[31:16]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_6 = _GEN_1 & 32'hffff; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_8 = {io_in1[15:0], 16'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_10 = _shin_T_8 & 32'hffff0000; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_11 = _shin_T_6 | _shin_T_10; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_2 = {{8'd0}, _shin_T_11[31:8]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_16 = _GEN_2 & 32'hff00ff; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_18 = {_shin_T_11[23:0], 8'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_20 = _shin_T_18 & 32'hff00ff00; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_21 = _shin_T_16 | _shin_T_20; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_3 = {{4'd0}, _shin_T_21[31:4]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_26 = _GEN_3 & 32'hf0f0f0f; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_28 = {_shin_T_21[27:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_30 = _shin_T_28 & 32'hf0f0f0f0; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_31 = _shin_T_26 | _shin_T_30; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_4 = {{2'd0}, _shin_T_31[31:2]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_36 = _GEN_4 & 32'h33333333; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_38 = {_shin_T_31[29:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_40 = _shin_T_38 & 32'hcccccccc; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_41 = _shin_T_36 | _shin_T_40; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_5 = {{1'd0}, _shin_T_41[31:1]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_46 = _GEN_5 & 32'h55555555; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_48 = {_shin_T_41[30:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_50 = _shin_T_48 & 32'haaaaaaaa; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_51 = _shin_T_46 | _shin_T_50; // @[Bitwise.scala 105:39]
  wire [31:0] shin = io_func == 5'h5 | io_func == 5'hb ? io_in1 : _shin_T_51; // @[ALU.scala 81:17]
  wire  _shout_r_T_4 = _in2_inv_T_2 & shin[31]; // @[ALU.scala 82:36]
  wire [32:0] _shout_r_T_6 = {_shout_r_T_4,shin}; // @[ALU.scala 82:57]
  wire [32:0] _shout_r_T_7 = $signed(_shout_r_T_6) >>> shamt; // @[ALU.scala 82:64]
  wire [31:0] shout_r = _shout_r_T_7[31:0]; // @[ALU.scala 82:73]
  wire [31:0] _GEN_6 = {{16'd0}, shout_r[31:16]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_3 = _GEN_6 & 32'hffff; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_5 = {shout_r[15:0], 16'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_7 = _shout_l_T_5 & 32'hffff0000; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_7 = {{8'd0}, _shout_l_T_8[31:8]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_13 = _GEN_7 & 32'hff00ff; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_15 = {_shout_l_T_8[23:0], 8'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_17 = _shout_l_T_15 & 32'hff00ff00; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_8 = {{4'd0}, _shout_l_T_18[31:4]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_23 = _GEN_8 & 32'hf0f0f0f; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_25 = {_shout_l_T_18[27:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_27 = _shout_l_T_25 & 32'hf0f0f0f0; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_9 = {{2'd0}, _shout_l_T_28[31:2]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_33 = _GEN_9 & 32'h33333333; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_35 = {_shout_l_T_28[29:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_37 = _shout_l_T_35 & 32'hcccccccc; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_10 = {{1'd0}, _shout_l_T_38[31:1]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_43 = _GEN_10 & 32'h55555555; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_45 = {_shout_l_T_38[30:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_47 = _shout_l_T_45 & 32'haaaaaaaa; // @[Bitwise.scala 105:80]
  wire [31:0] shout_l = _shout_l_T_43 | _shout_l_T_47; // @[Bitwise.scala 105:39]
  wire [31:0] _shout_T_3 = _shin_T_2 ? shout_r : 32'h0; // @[ALU.scala 84:18]
  wire [31:0] _shout_T_5 = io_func == 5'h1 ? shout_l : 32'h0; // @[ALU.scala 85:8]
  wire [31:0] shout = _shout_T_3 | _shout_T_5; // @[ALU.scala 84:82]
  wire [31:0] _logic_T_1 = io_in1 ^ io_in2; // @[ALU.scala 88:46]
  wire [31:0] _logic_T_3 = io_in1 | io_in2; // @[ALU.scala 89:35]
  wire [31:0] _logic_T_5 = io_in1 & io_in2; // @[ALU.scala 90:38]
  wire [31:0] _logic_T_6 = io_func == 5'h7 ? _logic_T_5 : 32'h0; // @[ALU.scala 90:10]
  wire [31:0] _logic_T_7 = io_func == 5'h6 ? _logic_T_3 : _logic_T_6; // @[ALU.scala 89:8]
  wire [31:0] logic_ = io_func == 5'h4 ? _logic_T_1 : _logic_T_7; // @[ALU.scala 88:18]
  wire  _shift_logic_cmp_T_2 = io_func >= 5'hc & _in2_inv_T_1; // @[ALU.scala 46:42]
  wire  _shift_logic_cmp_T_3 = _shift_logic_cmp_T_2 & slt; // @[ALU.scala 92:40]
  wire [31:0] _GEN_11 = {{31'd0}, _shift_logic_cmp_T_3}; // @[ALU.scala 92:47]
  wire [31:0] _shift_logic_cmp_T_4 = _GEN_11 | logic_; // @[ALU.scala 92:47]
  wire [31:0] shift_logic_cmp = _shift_logic_cmp_T_4 | shout; // @[ALU.scala 92:55]
  wire [31:0] out = io_func == 5'h0 | io_func == 5'ha ? adder_out : shift_logic_cmp; // @[ALU.scala 93:16]
  wire  _mul_in2_T = io_func == 5'h1a; // @[ALU.scala 97:26]
  wire  _mul_in2_T_2 = io_func == 5'h1a | io_func == 5'h1b; // @[ALU.scala 97:36]
  wire [31:0] mul_in2 = io_func == 5'h1a | io_func == 5'h1b ? io_in3 : io_in2; // @[ALU.scala 97:18]
  wire [63:0] in1_mul_in2_u = io_in1 * mul_in2; // @[ALU.scala 100:28]
  wire [31:0] _in1_mul_in2_T_1 = io_func == 5'h1a | io_func == 5'h1b ? io_in3 : io_in2; // @[ALU.scala 102:42]
  wire [63:0] in1_mul_in2 = $signed(io_in1) * $signed(_in1_mul_in2_T_1); // @[ALU.scala 102:32]
  wire [31:0] in1_mul_in2_l = in1_mul_in2[31:0]; // @[ALU.scala 103:32]
  wire [31:0] in1_mul_in2_h = in1_mul_in2[63:32]; // @[ALU.scala 104:32]
  wire [31:0] in1_mul_in2_hu = in1_mul_in2_u[63:32]; // @[ALU.scala 105:35]
  wire [32:0] _in1_mul_in2_hsu_T_1 = {1'b0,$signed(io_in1)}; // @[ALU.scala 106:40]
  wire [64:0] _in1_mul_in2_hsu_T_2 = $signed(_in1_mul_in2_T_1) * $signed(_in1_mul_in2_hsu_T_1); // @[ALU.scala 106:40]
  wire [63:0] _in1_mul_in2_hsu_T_4 = _in1_mul_in2_hsu_T_2[63:0]; // @[ALU.scala 106:40]
  wire [31:0] in1_mul_in2_hsu = _in1_mul_in2_hsu_T_4[63:32]; // @[ALU.scala 106:57]
  wire [31:0] _mul_out_T_3 = io_func == 5'h16 ? in1_mul_in2_hu : in1_mul_in2_hsu; // @[ALU.scala 109:20]
  wire [31:0] _mul_out_T_4 = io_func == 5'h15 ? in1_mul_in2_h : _mul_out_T_3; // @[ALU.scala 108:20]
  wire [31:0] mul_out = io_func == 5'h14 ? in1_mul_in2_l : _mul_out_T_4; // @[ALU.scala 107:20]
  wire [31:0] _in1_mul_in2_add_in3_T = in1_mul_in2[31:0]; // @[ALU.scala 111:44]
  wire [31:0] _in1_mul_in2_add_in3_T_1 = _mul_in2_T_2 ? io_in2 : io_in3; // @[ALU.scala 111:61]
  wire [31:0] in1_mul_in2_add_in3 = $signed(_in1_mul_in2_add_in3_T) + $signed(_in1_mul_in2_add_in3_T_1); // @[ALU.scala 111:68]
  wire [63:0] _GEN_12 = {{32{_in1_mul_in2_add_in3_T_1[31]}},_in1_mul_in2_add_in3_T_1}; // @[ALU.scala 112:52]
  wire [63:0] _minus_in1_mul_in2_add_in3_T_3 = $signed(_GEN_12) - $signed(in1_mul_in2); // @[ALU.scala 112:52]
  wire [31:0] minus_in1_mul_in2_add_in3 = _minus_in1_mul_in2_add_in3_T_3[31:0]; // @[ALU.scala 112:66]
  wire [31:0] mac_out = io_func == 5'h18 | _mul_in2_T ? in1_mul_in2_add_in3 : minus_in1_mul_in2_add_in3; // @[ALU.scala 116:20]
  wire  _minu_T = io_in1 > io_in2; // @[ALU.scala 119:22]
  wire [31:0] minu = io_in1 > io_in2 ? io_in2 : io_in1; // @[ALU.scala 119:15]
  wire [31:0] maxu = _minu_T ? io_in1 : io_in2; // @[ALU.scala 120:15]
  wire  _mins_T = $signed(io_in1) > $signed(io_in2); // @[ALU.scala 123:20]
  wire [31:0] mins = $signed(io_in1) > $signed(io_in2) ? $signed(io_in2) : $signed(io_in1); // @[ALU.scala 123:37]
  wire [31:0] maxs = _mins_T ? $signed(io_in1) : $signed(io_in2); // @[ALU.scala 124:37]
  wire [31:0] _minmaxout_T_3 = io_func == 5'h13 ? minu : maxu; // @[ALU.scala 127:22]
  wire [31:0] _minmaxout_T_4 = io_func == 5'h10 ? maxs : _minmaxout_T_3; // @[ALU.scala 126:22]
  wire [31:0] minmaxout = io_func == 5'h11 ? mins : _minmaxout_T_4; // @[ALU.scala 125:22]
  wire  _io_out_T_2 = io_func[4:2] == 3'h6; // @[ALU.scala 52:32]
  wire  _io_out_T_4 = io_func[4:2] == 3'h5; // @[ALU.scala 51:32]
  wire  _io_out_T_6 = io_func[4:2] == 3'h4; // @[ALU.scala 50:32]
  wire [31:0] _io_out_T_7 = _io_out_T_6 ? minmaxout : out; // @[ALU.scala 132:16]
  wire [31:0] _io_out_T_8 = _io_out_T_4 ? mul_out : _io_out_T_7; // @[ALU.scala 131:16]
  wire [31:0] _io_out_T_9 = _io_out_T_2 ? mac_out : _io_out_T_8; // @[ALU.scala 130:16]
  assign io_out = io_func == 5'h8 ? io_in2 : _io_out_T_9; // @[ALU.scala 129:16]
  assign io_cmp_out = io_func[0] ^ _io_cmp_out_T_4; // @[ALU.scala 77:38]
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_wb_wxd_rd,
  input         io_enq_bits_wxd,
  input  [4:0]  io_enq_bits_reg_idxw,
  input  [1:0]  io_enq_bits_warp_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_wb_wxd_rd,
  output        io_deq_bits_wxd,
  output [4:0]  io_deq_bits_reg_idxw,
  output [1:0]  io_deq_bits_warp_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_wb_wxd_rd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wxd_rd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wxd_rd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wxd_rd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wxd_rd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wxd_rd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wxd_rd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wxd_rd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wxd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wxd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wxd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wxd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wxd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wxd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wxd_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_reg_idxw [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_warp_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_warp_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_warp_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_wb_wxd_rd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wxd_rd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wxd_rd_io_deq_bits_MPORT_data = ram_wb_wxd_rd[ram_wb_wxd_rd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wxd_rd_MPORT_data = io_enq_bits_wb_wxd_rd;
  assign ram_wb_wxd_rd_MPORT_addr = 1'h0;
  assign ram_wb_wxd_rd_MPORT_mask = 1'h1;
  assign ram_wb_wxd_rd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wxd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wxd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wxd_io_deq_bits_MPORT_data = ram_wxd[ram_wxd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wxd_MPORT_data = io_enq_bits_wxd;
  assign ram_wxd_MPORT_addr = 1'h0;
  assign ram_wxd_MPORT_mask = 1'h1;
  assign ram_wxd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reg_idxw_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_reg_idxw_io_deq_bits_MPORT_data = ram_reg_idxw[ram_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_reg_idxw_MPORT_data = io_enq_bits_reg_idxw;
  assign ram_reg_idxw_MPORT_addr = 1'h0;
  assign ram_reg_idxw_MPORT_mask = 1'h1;
  assign ram_reg_idxw_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_warp_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_warp_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_warp_id_io_deq_bits_MPORT_data = ram_warp_id[ram_warp_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_warp_id_MPORT_data = io_enq_bits_warp_id;
  assign ram_warp_id_MPORT_addr = 1'h0;
  assign ram_warp_id_MPORT_mask = 1'h1;
  assign ram_warp_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_wb_wxd_rd = ram_wb_wxd_rd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wxd = ram_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_reg_idxw = ram_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_warp_id = ram_warp_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_wb_wxd_rd_MPORT_en & ram_wb_wxd_rd_MPORT_mask) begin
      ram_wb_wxd_rd[ram_wb_wxd_rd_MPORT_addr] <= ram_wb_wxd_rd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wxd_MPORT_en & ram_wxd_MPORT_mask) begin
      ram_wxd[ram_wxd_MPORT_addr] <= ram_wxd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_reg_idxw_MPORT_en & ram_reg_idxw_MPORT_mask) begin
      ram_reg_idxw[ram_reg_idxw_MPORT_addr] <= ram_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_warp_id_MPORT_en & ram_warp_id_MPORT_mask) begin
      ram_warp_id[ram_warp_id_MPORT_addr] <= ram_warp_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wxd_rd[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wxd[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_reg_idxw[initvar] = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_warp_id[initvar] = _RAND_3[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_wid,
  input         io_enq_bits_jump,
  input  [31:0] io_enq_bits_new_pc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_wid,
  output        io_deq_bits_jump,
  output [31:0] io_deq_bits_new_pc
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_jump [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_jump_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_jump_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_jump_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_new_pc [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_new_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_new_pc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wid_io_deq_bits_MPORT_data = ram_wid[ram_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wid_MPORT_data = io_enq_bits_wid;
  assign ram_wid_MPORT_addr = 1'h0;
  assign ram_wid_MPORT_mask = 1'h1;
  assign ram_wid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_jump_io_deq_bits_MPORT_en = 1'h1;
  assign ram_jump_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_jump_io_deq_bits_MPORT_data = ram_jump[ram_jump_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_jump_MPORT_data = io_enq_bits_jump;
  assign ram_jump_MPORT_addr = 1'h0;
  assign ram_jump_MPORT_mask = 1'h1;
  assign ram_jump_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_new_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_new_pc_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_new_pc_io_deq_bits_MPORT_data = ram_new_pc[ram_new_pc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_new_pc_MPORT_data = io_enq_bits_new_pc;
  assign ram_new_pc_MPORT_addr = 1'h0;
  assign ram_new_pc_MPORT_mask = 1'h1;
  assign ram_new_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_wid = ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_jump = ram_jump_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_new_pc = ram_new_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_wid_MPORT_en & ram_wid_MPORT_mask) begin
      ram_wid[ram_wid_MPORT_addr] <= ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_jump_MPORT_en & ram_jump_MPORT_mask) begin
      ram_jump[ram_jump_MPORT_addr] <= ram_jump_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_new_pc_MPORT_en & ram_new_pc_MPORT_mask) begin
      ram_new_pc[ram_new_pc_MPORT_addr] <= ram_new_pc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wid[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_jump[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_new_pc[initvar] = _RAND_2[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALUexe(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_in1,
  input  [31:0] io_in_bits_in2,
  input  [31:0] io_in_bits_in3,
  input  [1:0]  io_in_bits_ctrl_wid,
  input  [1:0]  io_in_bits_ctrl_branch,
  input  [5:0]  io_in_bits_ctrl_alu_fn,
  input  [4:0]  io_in_bits_ctrl_reg_idxw,
  input         io_in_bits_ctrl_wxd,
  output        io_out_valid,
  output [31:0] io_out_bits_wb_wxd_rd,
  output        io_out_bits_wxd,
  output [4:0]  io_out_bits_reg_idxw,
  output [1:0]  io_out_bits_warp_id,
  input         io_out2br_ready,
  output        io_out2br_valid,
  output [1:0]  io_out2br_bits_wid,
  output        io_out2br_bits_jump,
  output [31:0] io_out2br_bits_new_pc
);
  wire [4:0] alu_io_func; // @[execution.scala 19:17]
  wire [31:0] alu_io_in2; // @[execution.scala 19:17]
  wire [31:0] alu_io_in1; // @[execution.scala 19:17]
  wire [31:0] alu_io_in3; // @[execution.scala 19:17]
  wire [31:0] alu_io_out; // @[execution.scala 19:17]
  wire  alu_io_cmp_out; // @[execution.scala 19:17]
  wire  result_clock; // @[execution.scala 24:20]
  wire  result_reset; // @[execution.scala 24:20]
  wire  result_io_enq_ready; // @[execution.scala 24:20]
  wire  result_io_enq_valid; // @[execution.scala 24:20]
  wire [31:0] result_io_enq_bits_wb_wxd_rd; // @[execution.scala 24:20]
  wire  result_io_enq_bits_wxd; // @[execution.scala 24:20]
  wire [4:0] result_io_enq_bits_reg_idxw; // @[execution.scala 24:20]
  wire [1:0] result_io_enq_bits_warp_id; // @[execution.scala 24:20]
  wire  result_io_deq_ready; // @[execution.scala 24:20]
  wire  result_io_deq_valid; // @[execution.scala 24:20]
  wire [31:0] result_io_deq_bits_wb_wxd_rd; // @[execution.scala 24:20]
  wire  result_io_deq_bits_wxd; // @[execution.scala 24:20]
  wire [4:0] result_io_deq_bits_reg_idxw; // @[execution.scala 24:20]
  wire [1:0] result_io_deq_bits_warp_id; // @[execution.scala 24:20]
  wire  result_br_clock; // @[execution.scala 25:23]
  wire  result_br_reset; // @[execution.scala 25:23]
  wire  result_br_io_enq_ready; // @[execution.scala 25:23]
  wire  result_br_io_enq_valid; // @[execution.scala 25:23]
  wire [1:0] result_br_io_enq_bits_wid; // @[execution.scala 25:23]
  wire  result_br_io_enq_bits_jump; // @[execution.scala 25:23]
  wire [31:0] result_br_io_enq_bits_new_pc; // @[execution.scala 25:23]
  wire  result_br_io_deq_ready; // @[execution.scala 25:23]
  wire  result_br_io_deq_valid; // @[execution.scala 25:23]
  wire [1:0] result_br_io_deq_bits_wid; // @[execution.scala 25:23]
  wire  result_br_io_deq_bits_jump; // @[execution.scala 25:23]
  wire [31:0] result_br_io_deq_bits_new_pc; // @[execution.scala 25:23]
  wire  _io_in_ready_T = result_br_io_enq_ready & result_io_enq_ready; // @[execution.scala 34:71]
  wire  _io_in_ready_T_2 = 2'h1 == io_in_bits_ctrl_branch ? result_br_io_enq_ready : _io_in_ready_T; // @[Mux.scala 81:58]
  ScalarALU alu ( // @[execution.scala 19:17]
    .io_func(alu_io_func),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_in3(alu_io_in3),
    .io_out(alu_io_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  Queue_1 result ( // @[execution.scala 24:20]
    .clock(result_clock),
    .reset(result_reset),
    .io_enq_ready(result_io_enq_ready),
    .io_enq_valid(result_io_enq_valid),
    .io_enq_bits_wb_wxd_rd(result_io_enq_bits_wb_wxd_rd),
    .io_enq_bits_wxd(result_io_enq_bits_wxd),
    .io_enq_bits_reg_idxw(result_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_io_enq_bits_warp_id),
    .io_deq_ready(result_io_deq_ready),
    .io_deq_valid(result_io_deq_valid),
    .io_deq_bits_wb_wxd_rd(result_io_deq_bits_wb_wxd_rd),
    .io_deq_bits_wxd(result_io_deq_bits_wxd),
    .io_deq_bits_reg_idxw(result_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_io_deq_bits_warp_id)
  );
  Queue_2 result_br ( // @[execution.scala 25:23]
    .clock(result_br_clock),
    .reset(result_br_reset),
    .io_enq_ready(result_br_io_enq_ready),
    .io_enq_valid(result_br_io_enq_valid),
    .io_enq_bits_wid(result_br_io_enq_bits_wid),
    .io_enq_bits_jump(result_br_io_enq_bits_jump),
    .io_enq_bits_new_pc(result_br_io_enq_bits_new_pc),
    .io_deq_ready(result_br_io_deq_ready),
    .io_deq_valid(result_br_io_deq_valid),
    .io_deq_bits_wid(result_br_io_deq_bits_wid),
    .io_deq_bits_jump(result_br_io_deq_bits_jump),
    .io_deq_bits_new_pc(result_br_io_deq_bits_new_pc)
  );
  assign io_in_ready = 2'h0 == io_in_bits_ctrl_branch ? result_io_enq_ready : _io_in_ready_T_2; // @[Mux.scala 81:58]
  assign io_out_valid = result_io_deq_valid; // @[execution.scala 26:16]
  assign io_out_bits_wb_wxd_rd = result_io_deq_bits_wb_wxd_rd; // @[execution.scala 26:16]
  assign io_out_bits_wxd = result_io_deq_bits_wxd; // @[execution.scala 26:16]
  assign io_out_bits_reg_idxw = result_io_deq_bits_reg_idxw; // @[execution.scala 26:16]
  assign io_out_bits_warp_id = result_io_deq_bits_warp_id; // @[execution.scala 26:16]
  assign io_out2br_valid = result_br_io_deq_valid; // @[execution.scala 27:19]
  assign io_out2br_bits_wid = result_br_io_deq_bits_wid; // @[execution.scala 27:19]
  assign io_out2br_bits_jump = result_br_io_deq_bits_jump; // @[execution.scala 27:19]
  assign io_out2br_bits_new_pc = result_br_io_deq_bits_new_pc; // @[execution.scala 27:19]
  assign alu_io_func = io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 23:38]
  assign alu_io_in2 = io_in_bits_in2; // @[execution.scala 21:13]
  assign alu_io_in1 = io_in_bits_in1; // @[execution.scala 20:13]
  assign alu_io_in3 = io_in_bits_in3; // @[execution.scala 22:13]
  assign result_clock = clock;
  assign result_reset = reset;
  assign result_io_enq_valid = io_in_valid & io_in_bits_ctrl_wxd; // @[execution.scala 41:35]
  assign result_io_enq_bits_wb_wxd_rd = alu_io_out; // @[execution.scala 30:31]
  assign result_io_enq_bits_wxd = io_in_bits_ctrl_wxd; // @[execution.scala 32:25]
  assign result_io_enq_bits_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[execution.scala 31:30]
  assign result_io_enq_bits_warp_id = io_in_bits_ctrl_wid; // @[execution.scala 29:29]
  assign result_io_deq_ready = 1'h1; // @[execution.scala 26:16]
  assign result_br_clock = clock;
  assign result_br_reset = reset;
  assign result_br_io_enq_valid = io_in_valid & io_in_bits_ctrl_branch != 2'h0; // @[execution.scala 40:38]
  assign result_br_io_enq_bits_wid = io_in_bits_ctrl_wid; // @[execution.scala 36:28]
  assign result_br_io_enq_bits_jump = 2'h3 == io_in_bits_ctrl_branch | (2'h2 == io_in_bits_ctrl_branch | 2'h1 ==
    io_in_bits_ctrl_branch & alu_io_cmp_out); // @[Mux.scala 81:58]
  assign result_br_io_enq_bits_new_pc = io_in_bits_in3; // @[execution.scala 37:31]
  assign result_br_io_deq_ready = io_out2br_ready; // @[execution.scala 27:19]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_wb_wfd_rd_0,
  input  [31:0] io_enq_bits_wb_wfd_rd_1,
  input  [31:0] io_enq_bits_wb_wfd_rd_2,
  input  [31:0] io_enq_bits_wb_wfd_rd_3,
  input  [31:0] io_enq_bits_wb_wfd_rd_4,
  input  [31:0] io_enq_bits_wb_wfd_rd_5,
  input  [31:0] io_enq_bits_wb_wfd_rd_6,
  input  [31:0] io_enq_bits_wb_wfd_rd_7,
  input         io_enq_bits_wfd_mask_0,
  input         io_enq_bits_wfd_mask_1,
  input         io_enq_bits_wfd_mask_2,
  input         io_enq_bits_wfd_mask_3,
  input         io_enq_bits_wfd_mask_4,
  input         io_enq_bits_wfd_mask_5,
  input         io_enq_bits_wfd_mask_6,
  input         io_enq_bits_wfd_mask_7,
  input         io_enq_bits_wfd,
  input  [4:0]  io_enq_bits_reg_idxw,
  input  [1:0]  io_enq_bits_warp_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_wb_wfd_rd_0,
  output [31:0] io_deq_bits_wb_wfd_rd_1,
  output [31:0] io_deq_bits_wb_wfd_rd_2,
  output [31:0] io_deq_bits_wb_wfd_rd_3,
  output [31:0] io_deq_bits_wb_wfd_rd_4,
  output [31:0] io_deq_bits_wb_wfd_rd_5,
  output [31:0] io_deq_bits_wb_wfd_rd_6,
  output [31:0] io_deq_bits_wb_wfd_rd_7,
  output        io_deq_bits_wfd_mask_0,
  output        io_deq_bits_wfd_mask_1,
  output        io_deq_bits_wfd_mask_2,
  output        io_deq_bits_wfd_mask_3,
  output        io_deq_bits_wfd_mask_4,
  output        io_deq_bits_wfd_mask_5,
  output        io_deq_bits_wfd_mask_6,
  output        io_deq_bits_wfd_mask_7,
  output        io_deq_bits_wfd,
  output [4:0]  io_deq_bits_reg_idxw,
  output [1:0]  io_deq_bits_warp_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_wb_wfd_rd_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_wb_wfd_rd_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_wb_wfd_rd_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wb_wfd_rd_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd_mask_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_mask_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wfd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wfd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wfd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wfd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wfd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wfd_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_reg_idxw [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_reg_idxw_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_warp_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_warp_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_warp_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_warp_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_wb_wfd_rd_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_0_io_deq_bits_MPORT_data = ram_wb_wfd_rd_0[ram_wb_wfd_rd_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_0_MPORT_data = io_enq_bits_wb_wfd_rd_0;
  assign ram_wb_wfd_rd_0_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_0_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_1_io_deq_bits_MPORT_data = ram_wb_wfd_rd_1[ram_wb_wfd_rd_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_1_MPORT_data = io_enq_bits_wb_wfd_rd_1;
  assign ram_wb_wfd_rd_1_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_1_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_2_io_deq_bits_MPORT_data = ram_wb_wfd_rd_2[ram_wb_wfd_rd_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_2_MPORT_data = io_enq_bits_wb_wfd_rd_2;
  assign ram_wb_wfd_rd_2_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_2_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_3_io_deq_bits_MPORT_data = ram_wb_wfd_rd_3[ram_wb_wfd_rd_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_3_MPORT_data = io_enq_bits_wb_wfd_rd_3;
  assign ram_wb_wfd_rd_3_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_3_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_4_io_deq_bits_MPORT_data = ram_wb_wfd_rd_4[ram_wb_wfd_rd_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_4_MPORT_data = io_enq_bits_wb_wfd_rd_4;
  assign ram_wb_wfd_rd_4_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_4_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_5_io_deq_bits_MPORT_data = ram_wb_wfd_rd_5[ram_wb_wfd_rd_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_5_MPORT_data = io_enq_bits_wb_wfd_rd_5;
  assign ram_wb_wfd_rd_5_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_5_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_6_io_deq_bits_MPORT_data = ram_wb_wfd_rd_6[ram_wb_wfd_rd_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_6_MPORT_data = io_enq_bits_wb_wfd_rd_6;
  assign ram_wb_wfd_rd_6_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_6_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wb_wfd_rd_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wb_wfd_rd_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_7_io_deq_bits_MPORT_data = ram_wb_wfd_rd_7[ram_wb_wfd_rd_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wb_wfd_rd_7_MPORT_data = io_enq_bits_wb_wfd_rd_7;
  assign ram_wb_wfd_rd_7_MPORT_addr = 1'h0;
  assign ram_wb_wfd_rd_7_MPORT_mask = 1'h1;
  assign ram_wb_wfd_rd_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_0_io_deq_bits_MPORT_data = ram_wfd_mask_0[ram_wfd_mask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_0_MPORT_data = io_enq_bits_wfd_mask_0;
  assign ram_wfd_mask_0_MPORT_addr = 1'h0;
  assign ram_wfd_mask_0_MPORT_mask = 1'h1;
  assign ram_wfd_mask_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_1_io_deq_bits_MPORT_data = ram_wfd_mask_1[ram_wfd_mask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_1_MPORT_data = io_enq_bits_wfd_mask_1;
  assign ram_wfd_mask_1_MPORT_addr = 1'h0;
  assign ram_wfd_mask_1_MPORT_mask = 1'h1;
  assign ram_wfd_mask_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_2_io_deq_bits_MPORT_data = ram_wfd_mask_2[ram_wfd_mask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_2_MPORT_data = io_enq_bits_wfd_mask_2;
  assign ram_wfd_mask_2_MPORT_addr = 1'h0;
  assign ram_wfd_mask_2_MPORT_mask = 1'h1;
  assign ram_wfd_mask_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_3_io_deq_bits_MPORT_data = ram_wfd_mask_3[ram_wfd_mask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_3_MPORT_data = io_enq_bits_wfd_mask_3;
  assign ram_wfd_mask_3_MPORT_addr = 1'h0;
  assign ram_wfd_mask_3_MPORT_mask = 1'h1;
  assign ram_wfd_mask_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_4_io_deq_bits_MPORT_data = ram_wfd_mask_4[ram_wfd_mask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_4_MPORT_data = io_enq_bits_wfd_mask_4;
  assign ram_wfd_mask_4_MPORT_addr = 1'h0;
  assign ram_wfd_mask_4_MPORT_mask = 1'h1;
  assign ram_wfd_mask_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_5_io_deq_bits_MPORT_data = ram_wfd_mask_5[ram_wfd_mask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_5_MPORT_data = io_enq_bits_wfd_mask_5;
  assign ram_wfd_mask_5_MPORT_addr = 1'h0;
  assign ram_wfd_mask_5_MPORT_mask = 1'h1;
  assign ram_wfd_mask_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_6_io_deq_bits_MPORT_data = ram_wfd_mask_6[ram_wfd_mask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_6_MPORT_data = io_enq_bits_wfd_mask_6;
  assign ram_wfd_mask_6_MPORT_addr = 1'h0;
  assign ram_wfd_mask_6_MPORT_mask = 1'h1;
  assign ram_wfd_mask_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_mask_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_mask_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_mask_7_io_deq_bits_MPORT_data = ram_wfd_mask_7[ram_wfd_mask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_mask_7_MPORT_data = io_enq_bits_wfd_mask_7;
  assign ram_wfd_mask_7_MPORT_addr = 1'h0;
  assign ram_wfd_mask_7_MPORT_mask = 1'h1;
  assign ram_wfd_mask_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wfd_io_deq_bits_MPORT_data = ram_wfd[ram_wfd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wfd_MPORT_data = io_enq_bits_wfd;
  assign ram_wfd_MPORT_addr = 1'h0;
  assign ram_wfd_MPORT_mask = 1'h1;
  assign ram_wfd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reg_idxw_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_reg_idxw_io_deq_bits_MPORT_data = ram_reg_idxw[ram_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_reg_idxw_MPORT_data = io_enq_bits_reg_idxw;
  assign ram_reg_idxw_MPORT_addr = 1'h0;
  assign ram_reg_idxw_MPORT_mask = 1'h1;
  assign ram_reg_idxw_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_warp_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_warp_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_warp_id_io_deq_bits_MPORT_data = ram_warp_id[ram_warp_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_warp_id_MPORT_data = io_enq_bits_warp_id;
  assign ram_warp_id_MPORT_addr = 1'h0;
  assign ram_warp_id_MPORT_mask = 1'h1;
  assign ram_warp_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_wb_wfd_rd_0 = ram_wb_wfd_rd_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_1 = ram_wb_wfd_rd_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_2 = ram_wb_wfd_rd_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_3 = ram_wb_wfd_rd_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_4 = ram_wb_wfd_rd_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_5 = ram_wb_wfd_rd_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_6 = ram_wb_wfd_rd_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wb_wfd_rd_7 = ram_wb_wfd_rd_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_0 = ram_wfd_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_1 = ram_wfd_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_2 = ram_wfd_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_3 = ram_wfd_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_4 = ram_wfd_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_5 = ram_wfd_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_6 = ram_wfd_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd_mask_7 = ram_wfd_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wfd = ram_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_reg_idxw = ram_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_warp_id = ram_warp_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_wb_wfd_rd_0_MPORT_en & ram_wb_wfd_rd_0_MPORT_mask) begin
      ram_wb_wfd_rd_0[ram_wb_wfd_rd_0_MPORT_addr] <= ram_wb_wfd_rd_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_1_MPORT_en & ram_wb_wfd_rd_1_MPORT_mask) begin
      ram_wb_wfd_rd_1[ram_wb_wfd_rd_1_MPORT_addr] <= ram_wb_wfd_rd_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_2_MPORT_en & ram_wb_wfd_rd_2_MPORT_mask) begin
      ram_wb_wfd_rd_2[ram_wb_wfd_rd_2_MPORT_addr] <= ram_wb_wfd_rd_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_3_MPORT_en & ram_wb_wfd_rd_3_MPORT_mask) begin
      ram_wb_wfd_rd_3[ram_wb_wfd_rd_3_MPORT_addr] <= ram_wb_wfd_rd_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_4_MPORT_en & ram_wb_wfd_rd_4_MPORT_mask) begin
      ram_wb_wfd_rd_4[ram_wb_wfd_rd_4_MPORT_addr] <= ram_wb_wfd_rd_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_5_MPORT_en & ram_wb_wfd_rd_5_MPORT_mask) begin
      ram_wb_wfd_rd_5[ram_wb_wfd_rd_5_MPORT_addr] <= ram_wb_wfd_rd_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_6_MPORT_en & ram_wb_wfd_rd_6_MPORT_mask) begin
      ram_wb_wfd_rd_6[ram_wb_wfd_rd_6_MPORT_addr] <= ram_wb_wfd_rd_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wb_wfd_rd_7_MPORT_en & ram_wb_wfd_rd_7_MPORT_mask) begin
      ram_wb_wfd_rd_7[ram_wb_wfd_rd_7_MPORT_addr] <= ram_wb_wfd_rd_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_0_MPORT_en & ram_wfd_mask_0_MPORT_mask) begin
      ram_wfd_mask_0[ram_wfd_mask_0_MPORT_addr] <= ram_wfd_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_1_MPORT_en & ram_wfd_mask_1_MPORT_mask) begin
      ram_wfd_mask_1[ram_wfd_mask_1_MPORT_addr] <= ram_wfd_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_2_MPORT_en & ram_wfd_mask_2_MPORT_mask) begin
      ram_wfd_mask_2[ram_wfd_mask_2_MPORT_addr] <= ram_wfd_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_3_MPORT_en & ram_wfd_mask_3_MPORT_mask) begin
      ram_wfd_mask_3[ram_wfd_mask_3_MPORT_addr] <= ram_wfd_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_4_MPORT_en & ram_wfd_mask_4_MPORT_mask) begin
      ram_wfd_mask_4[ram_wfd_mask_4_MPORT_addr] <= ram_wfd_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_5_MPORT_en & ram_wfd_mask_5_MPORT_mask) begin
      ram_wfd_mask_5[ram_wfd_mask_5_MPORT_addr] <= ram_wfd_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_6_MPORT_en & ram_wfd_mask_6_MPORT_mask) begin
      ram_wfd_mask_6[ram_wfd_mask_6_MPORT_addr] <= ram_wfd_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_mask_7_MPORT_en & ram_wfd_mask_7_MPORT_mask) begin
      ram_wfd_mask_7[ram_wfd_mask_7_MPORT_addr] <= ram_wfd_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wfd_MPORT_en & ram_wfd_MPORT_mask) begin
      ram_wfd[ram_wfd_MPORT_addr] <= ram_wfd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_reg_idxw_MPORT_en & ram_reg_idxw_MPORT_mask) begin
      ram_reg_idxw[ram_reg_idxw_MPORT_addr] <= ram_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_warp_id_MPORT_en & ram_warp_id_MPORT_mask) begin
      ram_warp_id[ram_warp_id_MPORT_addr] <= ram_warp_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_0[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_1[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_2[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_3[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_4[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_5[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_6[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wb_wfd_rd_7[initvar] = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_0[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_1[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_2[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_3[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_4[initvar] = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_5[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_6[initvar] = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd_mask_7[initvar] = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wfd[initvar] = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_reg_idxw[initvar] = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_warp_id[initvar] = _RAND_18[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  maybe_full = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_if_mask,
  input  [1:0] io_enq_bits_wid,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_if_mask,
  output [1:0] io_deq_bits_wid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_if_mask [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_if_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_if_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_if_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_if_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_if_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_if_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_if_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_if_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_if_mask_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_if_mask_io_deq_bits_MPORT_data = ram_if_mask[ram_if_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_if_mask_MPORT_data = io_enq_bits_if_mask;
  assign ram_if_mask_MPORT_addr = 1'h0;
  assign ram_if_mask_MPORT_mask = 1'h1;
  assign ram_if_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wid_io_deq_bits_MPORT_data = ram_wid[ram_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wid_MPORT_data = io_enq_bits_wid;
  assign ram_wid_MPORT_addr = 1'h0;
  assign ram_wid_MPORT_mask = 1'h1;
  assign ram_wid_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_if_mask = ram_if_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_wid = ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_if_mask_MPORT_en & ram_if_mask_MPORT_mask) begin
      ram_if_mask[ram_if_mask_MPORT_addr] <= ram_if_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wid_MPORT_en & ram_wid_MPORT_mask) begin
      ram_wid[ram_wid_MPORT_addr] <= ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_if_mask[initvar] = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wid[initvar] = _RAND_1[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module vALUexe(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_in1_0,
  input  [31:0] io_in_bits_in1_1,
  input  [31:0] io_in_bits_in1_2,
  input  [31:0] io_in_bits_in1_3,
  input  [31:0] io_in_bits_in1_4,
  input  [31:0] io_in_bits_in1_5,
  input  [31:0] io_in_bits_in1_6,
  input  [31:0] io_in_bits_in1_7,
  input  [31:0] io_in_bits_in2_0,
  input  [31:0] io_in_bits_in2_1,
  input  [31:0] io_in_bits_in2_2,
  input  [31:0] io_in_bits_in2_3,
  input  [31:0] io_in_bits_in2_4,
  input  [31:0] io_in_bits_in2_5,
  input  [31:0] io_in_bits_in2_6,
  input  [31:0] io_in_bits_in2_7,
  input  [31:0] io_in_bits_in3_0,
  input  [31:0] io_in_bits_in3_1,
  input  [31:0] io_in_bits_in3_2,
  input  [31:0] io_in_bits_in3_3,
  input  [31:0] io_in_bits_in3_4,
  input  [31:0] io_in_bits_in3_5,
  input  [31:0] io_in_bits_in3_6,
  input  [31:0] io_in_bits_in3_7,
  input         io_in_bits_mask_0,
  input         io_in_bits_mask_1,
  input         io_in_bits_mask_2,
  input         io_in_bits_mask_3,
  input         io_in_bits_mask_4,
  input         io_in_bits_mask_5,
  input         io_in_bits_mask_6,
  input         io_in_bits_mask_7,
  input  [1:0]  io_in_bits_ctrl_wid,
  input         io_in_bits_ctrl_simt_stack,
  input         io_in_bits_ctrl_reverse,
  input  [5:0]  io_in_bits_ctrl_alu_fn,
  input  [4:0]  io_in_bits_ctrl_reg_idxw,
  input         io_in_bits_ctrl_wfd,
  input         io_in_bits_ctrl_readmask,
  input         io_in_bits_ctrl_writemask,
  output        io_out_valid,
  output [31:0] io_out_bits_wb_wfd_rd_0,
  output [31:0] io_out_bits_wb_wfd_rd_1,
  output [31:0] io_out_bits_wb_wfd_rd_2,
  output [31:0] io_out_bits_wb_wfd_rd_3,
  output [31:0] io_out_bits_wb_wfd_rd_4,
  output [31:0] io_out_bits_wb_wfd_rd_5,
  output [31:0] io_out_bits_wb_wfd_rd_6,
  output [31:0] io_out_bits_wb_wfd_rd_7,
  output        io_out_bits_wfd_mask_0,
  output        io_out_bits_wfd_mask_1,
  output        io_out_bits_wfd_mask_2,
  output        io_out_bits_wfd_mask_3,
  output        io_out_bits_wfd_mask_4,
  output        io_out_bits_wfd_mask_5,
  output        io_out_bits_wfd_mask_6,
  output        io_out_bits_wfd_mask_7,
  output        io_out_bits_wfd,
  output [4:0]  io_out_bits_reg_idxw,
  output [1:0]  io_out_bits_warp_id,
  input         io_out2simt_stack_ready,
  output        io_out2simt_stack_valid,
  output [7:0]  io_out2simt_stack_bits_if_mask,
  output [1:0]  io_out2simt_stack_bits_wid
);
  wire [4:0] ScalarALU_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_1_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_1_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_1_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_1_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_1_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_1_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_2_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_2_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_2_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_2_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_2_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_2_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_3_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_3_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_3_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_3_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_3_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_3_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_4_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_4_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_4_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_4_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_4_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_4_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_5_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_5_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_5_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_5_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_5_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_5_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_6_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_6_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_6_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_6_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_6_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_6_io_cmp_out; // @[execution.scala 50:47]
  wire [4:0] ScalarALU_7_io_func; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_7_io_in2; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_7_io_in1; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_7_io_in3; // @[execution.scala 50:47]
  wire [31:0] ScalarALU_7_io_out; // @[execution.scala 50:47]
  wire  ScalarALU_7_io_cmp_out; // @[execution.scala 50:47]
  wire  result_clock; // @[execution.scala 51:20]
  wire  result_reset; // @[execution.scala 51:20]
  wire  result_io_enq_ready; // @[execution.scala 51:20]
  wire  result_io_enq_valid; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_0; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_1; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_2; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_3; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_4; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_5; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_6; // @[execution.scala 51:20]
  wire [31:0] result_io_enq_bits_wb_wfd_rd_7; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_0; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_1; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_2; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_3; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_4; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_5; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_6; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd_mask_7; // @[execution.scala 51:20]
  wire  result_io_enq_bits_wfd; // @[execution.scala 51:20]
  wire [4:0] result_io_enq_bits_reg_idxw; // @[execution.scala 51:20]
  wire [1:0] result_io_enq_bits_warp_id; // @[execution.scala 51:20]
  wire  result_io_deq_ready; // @[execution.scala 51:20]
  wire  result_io_deq_valid; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_0; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_1; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_2; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_3; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_4; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_5; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_6; // @[execution.scala 51:20]
  wire [31:0] result_io_deq_bits_wb_wfd_rd_7; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_0; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_1; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_2; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_3; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_4; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_5; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_6; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd_mask_7; // @[execution.scala 51:20]
  wire  result_io_deq_bits_wfd; // @[execution.scala 51:20]
  wire [4:0] result_io_deq_bits_reg_idxw; // @[execution.scala 51:20]
  wire [1:0] result_io_deq_bits_warp_id; // @[execution.scala 51:20]
  wire  result2simt_clock; // @[execution.scala 52:25]
  wire  result2simt_reset; // @[execution.scala 52:25]
  wire  result2simt_io_enq_ready; // @[execution.scala 52:25]
  wire  result2simt_io_enq_valid; // @[execution.scala 52:25]
  wire [7:0] result2simt_io_enq_bits_if_mask; // @[execution.scala 52:25]
  wire [1:0] result2simt_io_enq_bits_wid; // @[execution.scala 52:25]
  wire  result2simt_io_deq_ready; // @[execution.scala 52:25]
  wire  result2simt_io_deq_valid; // @[execution.scala 52:25]
  wire [7:0] result2simt_io_deq_bits_if_mask; // @[execution.scala 52:25]
  wire [1:0] result2simt_io_deq_bits_wid; // @[execution.scala 52:25]
  wire [31:0] _GEN_0 = io_in_bits_ctrl_reverse ? io_in_bits_in2_0 : io_in_bits_in1_0; // @[execution.scala 54:15 59:34 60:17]
  wire  _T_2 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a; // @[execution.scala 63:48]
  wire  _T_3 = io_in_bits_ctrl_alu_fn == 6'h17; // @[execution.scala 63:110]
  wire  _T_5 = io_in_bits_ctrl_alu_fn == 6'h16; // @[execution.scala 63:147]
  wire  _T_7 = io_in_bits_ctrl_alu_fn == 6'h18; // @[execution.scala 63:183]
  wire [31:0] _alu_0_in1_T = ~io_in_bits_in1_0; // @[execution.scala 65:22]
  wire [4:0] _alu_0_func_T_2 = {4'h3,io_in_bits_ctrl_alu_fn[0]}; // @[Cat.scala 31:58]
  wire [4:0] _GEN_2 = _T_7 ? 5'h4 : _alu_0_func_T_2; // @[execution.scala 68:{49,61} 69:33]
  wire [31:0] alu_0_out = ScalarALU_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_0_T = ~alu_0_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_3 = _T_2 ? _alu_0_in1_T : _GEN_0; // @[execution.scala 64:89 65:19]
  wire [4:0] _GEN_4 = _T_2 ? _alu_0_func_T_2 : _GEN_2; // @[execution.scala 64:89 66:20]
  wire [31:0] _GEN_5 = _T_2 ? alu_0_out : _result_io_enq_bits_wb_wfd_rd_0_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_8 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_5 : alu_0_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_9 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h0 : _GEN_8; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_0_T_1 = io_in_bits_mask_0 ? io_in_bits_in1_0 : io_in_bits_in2_0; // @[execution.scala 77:43]
  wire [31:0] _GEN_10 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_0_T_1 : _GEN_9; // @[execution.scala 76:45 77:38]
  wire [31:0] _GEN_11 = io_in_bits_ctrl_reverse ? io_in_bits_in2_1 : io_in_bits_in1_1; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_1_in1_T = ~io_in_bits_in1_1; // @[execution.scala 65:22]
  wire [31:0] alu_1_out = ScalarALU_1_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_1_T = ~alu_1_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_14 = _T_2 ? _alu_1_in1_T : _GEN_11; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_16 = _T_2 ? alu_1_out : _result_io_enq_bits_wb_wfd_rd_1_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_19 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_16 : alu_1_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_20 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h1 : _GEN_19; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_1_T_1 = io_in_bits_mask_1 ? io_in_bits_in1_1 : io_in_bits_in2_1; // @[execution.scala 77:43]
  wire [31:0] _GEN_22 = io_in_bits_ctrl_reverse ? io_in_bits_in2_2 : io_in_bits_in1_2; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_2_in1_T = ~io_in_bits_in1_2; // @[execution.scala 65:22]
  wire [31:0] alu_2_out = ScalarALU_2_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_2_T = ~alu_2_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_25 = _T_2 ? _alu_2_in1_T : _GEN_22; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_27 = _T_2 ? alu_2_out : _result_io_enq_bits_wb_wfd_rd_2_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_30 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_27 : alu_2_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_31 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h2 : _GEN_30; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_2_T_1 = io_in_bits_mask_2 ? io_in_bits_in1_2 : io_in_bits_in2_2; // @[execution.scala 77:43]
  wire [31:0] _GEN_33 = io_in_bits_ctrl_reverse ? io_in_bits_in2_3 : io_in_bits_in1_3; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_3_in1_T = ~io_in_bits_in1_3; // @[execution.scala 65:22]
  wire [31:0] alu_3_out = ScalarALU_3_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_3_T = ~alu_3_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_36 = _T_2 ? _alu_3_in1_T : _GEN_33; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_38 = _T_2 ? alu_3_out : _result_io_enq_bits_wb_wfd_rd_3_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_41 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_38 : alu_3_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_42 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h3 : _GEN_41; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_3_T_1 = io_in_bits_mask_3 ? io_in_bits_in1_3 : io_in_bits_in2_3; // @[execution.scala 77:43]
  wire [31:0] _GEN_44 = io_in_bits_ctrl_reverse ? io_in_bits_in2_4 : io_in_bits_in1_4; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_4_in1_T = ~io_in_bits_in1_4; // @[execution.scala 65:22]
  wire [31:0] alu_4_out = ScalarALU_4_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_4_T = ~alu_4_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_47 = _T_2 ? _alu_4_in1_T : _GEN_44; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_49 = _T_2 ? alu_4_out : _result_io_enq_bits_wb_wfd_rd_4_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_52 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_49 : alu_4_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_53 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h4 : _GEN_52; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_4_T_1 = io_in_bits_mask_4 ? io_in_bits_in1_4 : io_in_bits_in2_4; // @[execution.scala 77:43]
  wire [31:0] _GEN_55 = io_in_bits_ctrl_reverse ? io_in_bits_in2_5 : io_in_bits_in1_5; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_5_in1_T = ~io_in_bits_in1_5; // @[execution.scala 65:22]
  wire [31:0] alu_5_out = ScalarALU_5_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_5_T = ~alu_5_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_58 = _T_2 ? _alu_5_in1_T : _GEN_55; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_60 = _T_2 ? alu_5_out : _result_io_enq_bits_wb_wfd_rd_5_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_63 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_60 : alu_5_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_64 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h5 : _GEN_63; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_5_T_1 = io_in_bits_mask_5 ? io_in_bits_in1_5 : io_in_bits_in2_5; // @[execution.scala 77:43]
  wire [31:0] _GEN_66 = io_in_bits_ctrl_reverse ? io_in_bits_in2_6 : io_in_bits_in1_6; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_6_in1_T = ~io_in_bits_in1_6; // @[execution.scala 65:22]
  wire [31:0] alu_6_out = ScalarALU_6_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_6_T = ~alu_6_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_69 = _T_2 ? _alu_6_in1_T : _GEN_66; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_71 = _T_2 ? alu_6_out : _result_io_enq_bits_wb_wfd_rd_6_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_74 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_71 : alu_6_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_75 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h6 : _GEN_74; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_6_T_1 = io_in_bits_mask_6 ? io_in_bits_in1_6 : io_in_bits_in2_6; // @[execution.scala 77:43]
  wire [31:0] _GEN_77 = io_in_bits_ctrl_reverse ? io_in_bits_in2_7 : io_in_bits_in1_7; // @[execution.scala 54:15 59:34 60:17]
  wire [31:0] _alu_7_in1_T = ~io_in_bits_in1_7; // @[execution.scala 65:22]
  wire [31:0] alu_7_out = ScalarALU_7_io_out; // @[execution.scala 50:{18,18}]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_7_T = ~alu_7_out; // @[execution.scala 70:43]
  wire [31:0] _GEN_80 = _T_2 ? _alu_7_in1_T : _GEN_77; // @[execution.scala 64:89 65:19]
  wire [31:0] _GEN_82 = _T_2 ? alu_7_out : _result_io_enq_bits_wb_wfd_rd_7_T; // @[execution.scala 58:36 64:89 70:40]
  wire [31:0] _GEN_85 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn == 6'h17
     | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_82 : alu_7_out; // @[execution.scala 63:197 58:36]
  wire [31:0] _GEN_86 = io_in_bits_ctrl_alu_fn == 6'h19 ? 32'h7 : _GEN_85; // @[execution.scala 73:42 74:38]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_7_T_1 = io_in_bits_mask_7 ? io_in_bits_in1_7 : io_in_bits_in2_7; // @[execution.scala 77:43]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_3 = io_in_bits_mask_0 & alu_0_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_5 = io_in_bits_mask_1 & alu_1_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_7 = io_in_bits_mask_2 & alu_2_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_9 = io_in_bits_mask_3 & alu_3_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_11 = io_in_bits_mask_4 & alu_4_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_13 = io_in_bits_mask_5 & alu_5_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_15 = io_in_bits_mask_6 & alu_6_out[0]; // @[execution.scala 82:118]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_17 = io_in_bits_mask_7 & alu_7_out[0]; // @[execution.scala 82:118]
  wire [7:0] _result_io_enq_bits_wb_wfd_rd_0_T_18 = {_result_io_enq_bits_wb_wfd_rd_0_T_17,
    _result_io_enq_bits_wb_wfd_rd_0_T_15,_result_io_enq_bits_wb_wfd_rd_0_T_13,_result_io_enq_bits_wb_wfd_rd_0_T_11,
    _result_io_enq_bits_wb_wfd_rd_0_T_9,_result_io_enq_bits_wb_wfd_rd_0_T_7,_result_io_enq_bits_wb_wfd_rd_0_T_5,
    _result_io_enq_bits_wb_wfd_rd_0_T_3}; // @[execution.scala 82:160]
  wire [31:0] _result_io_enq_bits_wb_wfd_rd_0_T_19 = io_in_bits_ctrl_readmask ? alu_0_out : {{24'd0},
    _result_io_enq_bits_wb_wfd_rd_0_T_18}; // @[execution.scala 82:41]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_22 = io_in_bits_mask_0 & ~alu_0_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_25 = io_in_bits_mask_1 & ~alu_1_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_28 = io_in_bits_mask_2 & ~alu_2_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_31 = io_in_bits_mask_3 & ~alu_3_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_34 = io_in_bits_mask_4 & ~alu_4_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_37 = io_in_bits_mask_5 & ~alu_5_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_40 = io_in_bits_mask_6 & ~alu_6_out[0]; // @[execution.scala 85:80]
  wire  _result_io_enq_bits_wb_wfd_rd_0_T_43 = io_in_bits_mask_7 & ~alu_7_out[0]; // @[execution.scala 85:80]
  wire [7:0] _result_io_enq_bits_wb_wfd_rd_0_T_44 = {_result_io_enq_bits_wb_wfd_rd_0_T_43,
    _result_io_enq_bits_wb_wfd_rd_0_T_40,_result_io_enq_bits_wb_wfd_rd_0_T_37,_result_io_enq_bits_wb_wfd_rd_0_T_34,
    _result_io_enq_bits_wb_wfd_rd_0_T_31,_result_io_enq_bits_wb_wfd_rd_0_T_28,_result_io_enq_bits_wb_wfd_rd_0_T_25,
    _result_io_enq_bits_wb_wfd_rd_0_T_22}; // @[execution.scala 85:127]
  wire [31:0] _GEN_88 = _T_3 | _T_5 | _T_7 ? {{24'd0}, _result_io_enq_bits_wb_wfd_rd_0_T_44} :
    _result_io_enq_bits_wb_wfd_rd_0_T_19; // @[execution.scala 84:120 82:36 85:38]
  wire  alu_1_cmp_out = ScalarALU_1_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_0_cmp_out = ScalarALU_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_3_cmp_out = ScalarALU_3_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_2_cmp_out = ScalarALU_2_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_5_cmp_out = ScalarALU_5_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_4_cmp_out = ScalarALU_4_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_7_cmp_out = ScalarALU_7_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire  alu_6_cmp_out = ScalarALU_6_io_cmp_out; // @[execution.scala 50:{18,18}]
  wire [7:0] _result2simt_io_enq_bits_if_mask_T = {alu_7_cmp_out,alu_6_cmp_out,alu_5_cmp_out,alu_4_cmp_out,alu_3_cmp_out
    ,alu_2_cmp_out,alu_1_cmp_out,alu_0_cmp_out}; // @[execution.scala 96:72]
  ScalarALU ScalarALU ( // @[execution.scala 50:47]
    .io_func(ScalarALU_io_func),
    .io_in2(ScalarALU_io_in2),
    .io_in1(ScalarALU_io_in1),
    .io_in3(ScalarALU_io_in3),
    .io_out(ScalarALU_io_out),
    .io_cmp_out(ScalarALU_io_cmp_out)
  );
  ScalarALU ScalarALU_1 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_1_io_func),
    .io_in2(ScalarALU_1_io_in2),
    .io_in1(ScalarALU_1_io_in1),
    .io_in3(ScalarALU_1_io_in3),
    .io_out(ScalarALU_1_io_out),
    .io_cmp_out(ScalarALU_1_io_cmp_out)
  );
  ScalarALU ScalarALU_2 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_2_io_func),
    .io_in2(ScalarALU_2_io_in2),
    .io_in1(ScalarALU_2_io_in1),
    .io_in3(ScalarALU_2_io_in3),
    .io_out(ScalarALU_2_io_out),
    .io_cmp_out(ScalarALU_2_io_cmp_out)
  );
  ScalarALU ScalarALU_3 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_3_io_func),
    .io_in2(ScalarALU_3_io_in2),
    .io_in1(ScalarALU_3_io_in1),
    .io_in3(ScalarALU_3_io_in3),
    .io_out(ScalarALU_3_io_out),
    .io_cmp_out(ScalarALU_3_io_cmp_out)
  );
  ScalarALU ScalarALU_4 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_4_io_func),
    .io_in2(ScalarALU_4_io_in2),
    .io_in1(ScalarALU_4_io_in1),
    .io_in3(ScalarALU_4_io_in3),
    .io_out(ScalarALU_4_io_out),
    .io_cmp_out(ScalarALU_4_io_cmp_out)
  );
  ScalarALU ScalarALU_5 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_5_io_func),
    .io_in2(ScalarALU_5_io_in2),
    .io_in1(ScalarALU_5_io_in1),
    .io_in3(ScalarALU_5_io_in3),
    .io_out(ScalarALU_5_io_out),
    .io_cmp_out(ScalarALU_5_io_cmp_out)
  );
  ScalarALU ScalarALU_6 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_6_io_func),
    .io_in2(ScalarALU_6_io_in2),
    .io_in1(ScalarALU_6_io_in1),
    .io_in3(ScalarALU_6_io_in3),
    .io_out(ScalarALU_6_io_out),
    .io_cmp_out(ScalarALU_6_io_cmp_out)
  );
  ScalarALU ScalarALU_7 ( // @[execution.scala 50:47]
    .io_func(ScalarALU_7_io_func),
    .io_in2(ScalarALU_7_io_in2),
    .io_in1(ScalarALU_7_io_in1),
    .io_in3(ScalarALU_7_io_in3),
    .io_out(ScalarALU_7_io_out),
    .io_cmp_out(ScalarALU_7_io_cmp_out)
  );
  Queue_3 result ( // @[execution.scala 51:20]
    .clock(result_clock),
    .reset(result_reset),
    .io_enq_ready(result_io_enq_ready),
    .io_enq_valid(result_io_enq_valid),
    .io_enq_bits_wb_wfd_rd_0(result_io_enq_bits_wb_wfd_rd_0),
    .io_enq_bits_wb_wfd_rd_1(result_io_enq_bits_wb_wfd_rd_1),
    .io_enq_bits_wb_wfd_rd_2(result_io_enq_bits_wb_wfd_rd_2),
    .io_enq_bits_wb_wfd_rd_3(result_io_enq_bits_wb_wfd_rd_3),
    .io_enq_bits_wb_wfd_rd_4(result_io_enq_bits_wb_wfd_rd_4),
    .io_enq_bits_wb_wfd_rd_5(result_io_enq_bits_wb_wfd_rd_5),
    .io_enq_bits_wb_wfd_rd_6(result_io_enq_bits_wb_wfd_rd_6),
    .io_enq_bits_wb_wfd_rd_7(result_io_enq_bits_wb_wfd_rd_7),
    .io_enq_bits_wfd_mask_0(result_io_enq_bits_wfd_mask_0),
    .io_enq_bits_wfd_mask_1(result_io_enq_bits_wfd_mask_1),
    .io_enq_bits_wfd_mask_2(result_io_enq_bits_wfd_mask_2),
    .io_enq_bits_wfd_mask_3(result_io_enq_bits_wfd_mask_3),
    .io_enq_bits_wfd_mask_4(result_io_enq_bits_wfd_mask_4),
    .io_enq_bits_wfd_mask_5(result_io_enq_bits_wfd_mask_5),
    .io_enq_bits_wfd_mask_6(result_io_enq_bits_wfd_mask_6),
    .io_enq_bits_wfd_mask_7(result_io_enq_bits_wfd_mask_7),
    .io_enq_bits_wfd(result_io_enq_bits_wfd),
    .io_enq_bits_reg_idxw(result_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_io_enq_bits_warp_id),
    .io_deq_ready(result_io_deq_ready),
    .io_deq_valid(result_io_deq_valid),
    .io_deq_bits_wb_wfd_rd_0(result_io_deq_bits_wb_wfd_rd_0),
    .io_deq_bits_wb_wfd_rd_1(result_io_deq_bits_wb_wfd_rd_1),
    .io_deq_bits_wb_wfd_rd_2(result_io_deq_bits_wb_wfd_rd_2),
    .io_deq_bits_wb_wfd_rd_3(result_io_deq_bits_wb_wfd_rd_3),
    .io_deq_bits_wb_wfd_rd_4(result_io_deq_bits_wb_wfd_rd_4),
    .io_deq_bits_wb_wfd_rd_5(result_io_deq_bits_wb_wfd_rd_5),
    .io_deq_bits_wb_wfd_rd_6(result_io_deq_bits_wb_wfd_rd_6),
    .io_deq_bits_wb_wfd_rd_7(result_io_deq_bits_wb_wfd_rd_7),
    .io_deq_bits_wfd_mask_0(result_io_deq_bits_wfd_mask_0),
    .io_deq_bits_wfd_mask_1(result_io_deq_bits_wfd_mask_1),
    .io_deq_bits_wfd_mask_2(result_io_deq_bits_wfd_mask_2),
    .io_deq_bits_wfd_mask_3(result_io_deq_bits_wfd_mask_3),
    .io_deq_bits_wfd_mask_4(result_io_deq_bits_wfd_mask_4),
    .io_deq_bits_wfd_mask_5(result_io_deq_bits_wfd_mask_5),
    .io_deq_bits_wfd_mask_6(result_io_deq_bits_wfd_mask_6),
    .io_deq_bits_wfd_mask_7(result_io_deq_bits_wfd_mask_7),
    .io_deq_bits_wfd(result_io_deq_bits_wfd),
    .io_deq_bits_reg_idxw(result_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_io_deq_bits_warp_id)
  );
  Queue_4 result2simt ( // @[execution.scala 52:25]
    .clock(result2simt_clock),
    .reset(result2simt_reset),
    .io_enq_ready(result2simt_io_enq_ready),
    .io_enq_valid(result2simt_io_enq_valid),
    .io_enq_bits_if_mask(result2simt_io_enq_bits_if_mask),
    .io_enq_bits_wid(result2simt_io_enq_bits_wid),
    .io_deq_ready(result2simt_io_deq_ready),
    .io_deq_valid(result2simt_io_deq_valid),
    .io_deq_bits_if_mask(result2simt_io_deq_bits_if_mask),
    .io_deq_bits_wid(result2simt_io_deq_bits_wid)
  );
  assign io_in_ready = io_in_bits_ctrl_simt_stack ? result2simt_io_enq_ready : result_io_enq_ready; // @[execution.scala 99:19]
  assign io_out_valid = result_io_deq_valid; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_0 = result_io_deq_bits_wb_wfd_rd_0; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_1 = result_io_deq_bits_wb_wfd_rd_1; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_2 = result_io_deq_bits_wb_wfd_rd_2; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_3 = result_io_deq_bits_wb_wfd_rd_3; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_4 = result_io_deq_bits_wb_wfd_rd_4; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_5 = result_io_deq_bits_wb_wfd_rd_5; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_6 = result_io_deq_bits_wb_wfd_rd_6; // @[execution.scala 100:9]
  assign io_out_bits_wb_wfd_rd_7 = result_io_deq_bits_wb_wfd_rd_7; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_0 = result_io_deq_bits_wfd_mask_0; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_1 = result_io_deq_bits_wfd_mask_1; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_2 = result_io_deq_bits_wfd_mask_2; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_3 = result_io_deq_bits_wfd_mask_3; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_4 = result_io_deq_bits_wfd_mask_4; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_5 = result_io_deq_bits_wfd_mask_5; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_6 = result_io_deq_bits_wfd_mask_6; // @[execution.scala 100:9]
  assign io_out_bits_wfd_mask_7 = result_io_deq_bits_wfd_mask_7; // @[execution.scala 100:9]
  assign io_out_bits_wfd = result_io_deq_bits_wfd; // @[execution.scala 100:9]
  assign io_out_bits_reg_idxw = result_io_deq_bits_reg_idxw; // @[execution.scala 100:9]
  assign io_out_bits_warp_id = result_io_deq_bits_warp_id; // @[execution.scala 100:9]
  assign io_out2simt_stack_valid = result2simt_io_deq_valid; // @[execution.scala 101:20]
  assign io_out2simt_stack_bits_if_mask = result2simt_io_deq_bits_if_mask; // @[execution.scala 101:20]
  assign io_out2simt_stack_bits_wid = result2simt_io_deq_bits_wid; // @[execution.scala 101:20]
  assign ScalarALU_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 : io_in_bits_ctrl_alu_fn[4:0]
    ; // @[execution.scala 57:16 63:197]
  assign ScalarALU_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_0 : io_in_bits_in2_0; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_3 : _GEN_0; // @[execution.scala 63:197]
  assign ScalarALU_io_in3 = io_in_bits_in3_0; // @[execution.scala 50:18 56:15]
  assign ScalarALU_1_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_1_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_1 : io_in_bits_in2_1; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_1_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_14 : _GEN_11; // @[execution.scala 63:197]
  assign ScalarALU_1_io_in3 = io_in_bits_in3_1; // @[execution.scala 50:18 56:15]
  assign ScalarALU_2_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_2_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_2 : io_in_bits_in2_2; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_2_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_25 : _GEN_22; // @[execution.scala 63:197]
  assign ScalarALU_2_io_in3 = io_in_bits_in3_2; // @[execution.scala 50:18 56:15]
  assign ScalarALU_3_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_3_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_3 : io_in_bits_in2_3; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_3_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_36 : _GEN_33; // @[execution.scala 63:197]
  assign ScalarALU_3_io_in3 = io_in_bits_in3_3; // @[execution.scala 50:18 56:15]
  assign ScalarALU_4_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_4_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_4 : io_in_bits_in2_4; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_4_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_47 : _GEN_44; // @[execution.scala 63:197]
  assign ScalarALU_4_io_in3 = io_in_bits_in3_4; // @[execution.scala 50:18 56:15]
  assign ScalarALU_5_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_5_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_5 : io_in_bits_in2_5; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_5_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_58 : _GEN_55; // @[execution.scala 63:197]
  assign ScalarALU_5_io_in3 = io_in_bits_in3_5; // @[execution.scala 50:18 56:15]
  assign ScalarALU_6_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_6_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_6 : io_in_bits_in2_6; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_6_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_69 : _GEN_66; // @[execution.scala 63:197]
  assign ScalarALU_6_io_in3 = io_in_bits_in3_6; // @[execution.scala 50:18 56:15]
  assign ScalarALU_7_io_func = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a |
    io_in_bits_ctrl_alu_fn == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_4 :
    io_in_bits_ctrl_alu_fn[4:0]; // @[execution.scala 57:16 63:197]
  assign ScalarALU_7_io_in2 = io_in_bits_ctrl_reverse ? io_in_bits_in1_7 : io_in_bits_in2_7; // @[execution.scala 55:15 59:34 61:17]
  assign ScalarALU_7_io_in1 = io_in_bits_ctrl_alu_fn == 6'h1b | io_in_bits_ctrl_alu_fn == 6'h1a | io_in_bits_ctrl_alu_fn
     == 6'h17 | io_in_bits_ctrl_alu_fn == 6'h16 | io_in_bits_ctrl_alu_fn == 6'h18 ? _GEN_80 : _GEN_77; // @[execution.scala 63:197]
  assign ScalarALU_7_io_in3 = io_in_bits_in3_7; // @[execution.scala 50:18 56:15]
  assign result_clock = clock;
  assign result_reset = reset;
  assign result_io_enq_valid = io_in_valid & io_in_bits_ctrl_wfd & ~io_in_bits_ctrl_simt_stack; // @[execution.scala 93:55]
  assign result_io_enq_bits_wb_wfd_rd_0 = io_in_bits_ctrl_writemask ? _GEN_88 : _GEN_10; // @[execution.scala 81:34]
  assign result_io_enq_bits_wb_wfd_rd_1 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_1_T_1 :
    _GEN_20; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wb_wfd_rd_2 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_2_T_1 :
    _GEN_31; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wb_wfd_rd_3 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_3_T_1 :
    _GEN_42; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wb_wfd_rd_4 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_4_T_1 :
    _GEN_53; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wb_wfd_rd_5 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_5_T_1 :
    _GEN_64; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wb_wfd_rd_6 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_6_T_1 :
    _GEN_75; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wb_wfd_rd_7 = io_in_bits_ctrl_alu_fn == 6'h13 ? _result_io_enq_bits_wb_wfd_rd_7_T_1 :
    _GEN_86; // @[execution.scala 76:45 77:38]
  assign result_io_enq_bits_wfd_mask_0 = io_in_bits_mask_0; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_1 = io_in_bits_mask_1; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_2 = io_in_bits_mask_2; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_3 = io_in_bits_mask_3; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_4 = io_in_bits_mask_4; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_5 = io_in_bits_mask_5; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_6 = io_in_bits_mask_6; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd_mask_7 = io_in_bits_mask_7; // @[execution.scala 92:30]
  assign result_io_enq_bits_wfd = io_in_bits_ctrl_wfd; // @[execution.scala 91:25]
  assign result_io_enq_bits_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[execution.scala 90:30]
  assign result_io_enq_bits_warp_id = io_in_bits_ctrl_wid; // @[execution.scala 89:29]
  assign result_io_deq_ready = 1'h1; // @[execution.scala 100:9]
  assign result2simt_clock = clock;
  assign result2simt_reset = reset;
  assign result2simt_io_enq_valid = io_in_valid & io_in_bits_ctrl_simt_stack; // @[execution.scala 97:40]
  assign result2simt_io_enq_bits_if_mask = ~_result2simt_io_enq_bits_if_mask_T; // @[execution.scala 96:37]
  assign result2simt_io_enq_bits_wid = io_in_bits_ctrl_wid; // @[execution.scala 95:30]
  assign result2simt_io_deq_ready = io_out2simt_stack_ready; // @[execution.scala 101:20]
endmodule
module Classify(
  input  [31:0] io_in,
  output        io_isNegInf,
  output        io_isNegNormal,
  output        io_isNegSubnormal,
  output        io_isNegZero,
  output        io_isPosZero,
  output        io_isPosSubnormal,
  output        io_isPosNormal,
  output        io_isPosInf,
  output        io_isSNaN,
  output        io_isQNaN,
  output        io_isNaN,
  output        io_isInf,
  output        io_isInfOrNaN,
  output        io_isSubnormal,
  output        io_isZero,
  output        io_isSubnormalOrZero
);
  wire [22:0] flpt_frac = io_in[22:0]; // @[Classify.scala 27:28]
  wire [7:0] flpt_exp = io_in[30:23]; // @[Classify.scala 27:28]
  wire  flpt_sign = io_in[31]; // @[Classify.scala 27:28]
  wire  isSubnormalOrZero = flpt_exp == 8'h0; // @[Classify.scala 30:31]
  wire  fracIsZero = flpt_frac == 23'h0; // @[Classify.scala 31:25]
  wire [7:0] _isInfOrNaN_T = ~flpt_exp; // @[Classify.scala 32:21]
  wire  isInfOrNaN = _isInfOrNaN_T == 8'h0; // @[Classify.scala 32:36]
  wire  _io_isNegNormal_T = ~isSubnormalOrZero; // @[Classify.scala 35:29]
  wire  _io_isNegNormal_T_2 = ~isInfOrNaN; // @[Classify.scala 35:51]
  wire  _io_isPosInf_T = ~flpt_sign; // @[Classify.scala 39:18]
  wire  _io_isNaN_T = ~fracIsZero; // @[Classify.scala 47:29]
  assign io_isNegInf = flpt_sign & io_isInf; // @[Classify.scala 34:23]
  assign io_isNegNormal = flpt_sign & ~isSubnormalOrZero & ~isInfOrNaN; // @[Classify.scala 35:48]
  assign io_isNegSubnormal = flpt_sign & io_isSubnormal; // @[Classify.scala 36:29]
  assign io_isNegZero = flpt_sign & io_isZero; // @[Classify.scala 37:24]
  assign io_isPosZero = _io_isPosInf_T & io_isZero; // @[Classify.scala 42:25]
  assign io_isPosSubnormal = _io_isPosInf_T & io_isSubnormal; // @[Classify.scala 41:30]
  assign io_isPosNormal = _io_isPosInf_T & _io_isNegNormal_T & _io_isNegNormal_T_2; // @[Classify.scala 40:49]
  assign io_isPosInf = ~flpt_sign & io_isInf; // @[Classify.scala 39:24]
  assign io_isSNaN = io_isNaN & ~flpt_frac[22]; // @[Classify.scala 44:25]
  assign io_isQNaN = io_isNaN & flpt_frac[22]; // @[Classify.scala 45:25]
  assign io_isNaN = isInfOrNaN & ~fracIsZero; // @[Classify.scala 47:26]
  assign io_isInf = isInfOrNaN & fracIsZero; // @[Classify.scala 48:26]
  assign io_isInfOrNaN = _isInfOrNaN_T == 8'h0; // @[Classify.scala 32:36]
  assign io_isSubnormal = isSubnormalOrZero & _io_isNaN_T; // @[Classify.scala 51:39]
  assign io_isZero = isSubnormalOrZero & fracIsZero; // @[Classify.scala 52:34]
  assign io_isSubnormalOrZero = flpt_exp == 8'h0; // @[Classify.scala 30:31]
endmodule
module ArrayMultiplier(
  input  [24:0] io_a,
  input  [24:0] io_b,
  output [49:0] io_sum
);
  assign io_sum = io_a * io_b; // @[FPU.scala 60:24]
endmodule
module RoundingUnit(
  input  [2:0]  io_in_rm,
  input  [23:0] io_in_frac,
  input         io_in_sign,
  input         io_in_guard,
  input         io_in_round,
  input         io_in_sticky,
  output [23:0] io_out_fracRounded,
  output        io_out_fracCout
);
  wire  inexact = io_in_guard | io_in_round | io_in_sticky; // @[FPU.scala 36:43]
  wire  lsb = io_in_frac[0]; // @[FPU.scala 37:23]
  wire  _roundUp_T_2 = io_in_guard & (io_in_round | io_in_sticky | lsb); // @[FPU.scala 39:25]
  wire  _roundUp_T_4 = inexact & ~io_in_sign; // @[FPU.scala 41:21]
  wire  _roundUp_T_5 = inexact & io_in_sign; // @[FPU.scala 42:21]
  wire  _roundUp_T_9 = 3'h1 == io_in_rm ? 1'h0 : 3'h0 == io_in_rm & _roundUp_T_2; // @[Mux.scala 81:58]
  wire  _roundUp_T_11 = 3'h3 == io_in_rm ? _roundUp_T_4 : _roundUp_T_9; // @[Mux.scala 81:58]
  wire  _roundUp_T_13 = 3'h2 == io_in_rm ? _roundUp_T_5 : _roundUp_T_11; // @[Mux.scala 81:58]
  wire  roundUp = 3'h4 == io_in_rm ? io_in_guard : _roundUp_T_13; // @[Mux.scala 81:58]
  wire [24:0] fracRoundUp = io_in_frac + 24'h1; // @[FPU.scala 45:32]
  wire  cout = fracRoundUp[24]; // @[FPU.scala 46:25]
  assign io_out_fracRounded = roundUp ? fracRoundUp[23:0] : io_in_frac; // @[FPU.scala 47:24]
  assign io_out_fracCout = cout & roundUp; // @[FPU.scala 50:27]
endmodule
module FPU_FMA(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_op,
  input  [31:0] io_in_bits_a,
  input  [31:0] io_in_bits_b,
  input  [31:0] io_in_bits_c,
  input  [2:0]  io_in_bits_rm,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [95:0] _RAND_26;
  reg [95:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] Classify_io_in; // @[FPU.scala 99:38]
  wire  Classify_io_isNegInf; // @[FPU.scala 99:38]
  wire  Classify_io_isNegNormal; // @[FPU.scala 99:38]
  wire  Classify_io_isNegSubnormal; // @[FPU.scala 99:38]
  wire  Classify_io_isNegZero; // @[FPU.scala 99:38]
  wire  Classify_io_isPosZero; // @[FPU.scala 99:38]
  wire  Classify_io_isPosSubnormal; // @[FPU.scala 99:38]
  wire  Classify_io_isPosNormal; // @[FPU.scala 99:38]
  wire  Classify_io_isPosInf; // @[FPU.scala 99:38]
  wire  Classify_io_isSNaN; // @[FPU.scala 99:38]
  wire  Classify_io_isQNaN; // @[FPU.scala 99:38]
  wire  Classify_io_isNaN; // @[FPU.scala 99:38]
  wire  Classify_io_isInf; // @[FPU.scala 99:38]
  wire  Classify_io_isInfOrNaN; // @[FPU.scala 99:38]
  wire  Classify_io_isSubnormal; // @[FPU.scala 99:38]
  wire  Classify_io_isZero; // @[FPU.scala 99:38]
  wire  Classify_io_isSubnormalOrZero; // @[FPU.scala 99:38]
  wire [31:0] Classify_1_io_in; // @[FPU.scala 99:38]
  wire  Classify_1_io_isNegInf; // @[FPU.scala 99:38]
  wire  Classify_1_io_isNegNormal; // @[FPU.scala 99:38]
  wire  Classify_1_io_isNegSubnormal; // @[FPU.scala 99:38]
  wire  Classify_1_io_isNegZero; // @[FPU.scala 99:38]
  wire  Classify_1_io_isPosZero; // @[FPU.scala 99:38]
  wire  Classify_1_io_isPosSubnormal; // @[FPU.scala 99:38]
  wire  Classify_1_io_isPosNormal; // @[FPU.scala 99:38]
  wire  Classify_1_io_isPosInf; // @[FPU.scala 99:38]
  wire  Classify_1_io_isSNaN; // @[FPU.scala 99:38]
  wire  Classify_1_io_isQNaN; // @[FPU.scala 99:38]
  wire  Classify_1_io_isNaN; // @[FPU.scala 99:38]
  wire  Classify_1_io_isInf; // @[FPU.scala 99:38]
  wire  Classify_1_io_isInfOrNaN; // @[FPU.scala 99:38]
  wire  Classify_1_io_isSubnormal; // @[FPU.scala 99:38]
  wire  Classify_1_io_isZero; // @[FPU.scala 99:38]
  wire  Classify_1_io_isSubnormalOrZero; // @[FPU.scala 99:38]
  wire [31:0] Classify_2_io_in; // @[FPU.scala 99:38]
  wire  Classify_2_io_isNegInf; // @[FPU.scala 99:38]
  wire  Classify_2_io_isNegNormal; // @[FPU.scala 99:38]
  wire  Classify_2_io_isNegSubnormal; // @[FPU.scala 99:38]
  wire  Classify_2_io_isNegZero; // @[FPU.scala 99:38]
  wire  Classify_2_io_isPosZero; // @[FPU.scala 99:38]
  wire  Classify_2_io_isPosSubnormal; // @[FPU.scala 99:38]
  wire  Classify_2_io_isPosNormal; // @[FPU.scala 99:38]
  wire  Classify_2_io_isPosInf; // @[FPU.scala 99:38]
  wire  Classify_2_io_isSNaN; // @[FPU.scala 99:38]
  wire  Classify_2_io_isQNaN; // @[FPU.scala 99:38]
  wire  Classify_2_io_isNaN; // @[FPU.scala 99:38]
  wire  Classify_2_io_isInf; // @[FPU.scala 99:38]
  wire  Classify_2_io_isInfOrNaN; // @[FPU.scala 99:38]
  wire  Classify_2_io_isSubnormal; // @[FPU.scala 99:38]
  wire  Classify_2_io_isZero; // @[FPU.scala 99:38]
  wire  Classify_2_io_isSubnormalOrZero; // @[FPU.scala 99:38]
  wire [24:0] mult_io_a; // @[FPU.scala 155:20]
  wire [24:0] mult_io_b; // @[FPU.scala 155:20]
  wire [49:0] mult_io_sum; // @[FPU.scala 155:20]
  wire [2:0] rounding_io_in_rm; // @[FPU.scala 274:24]
  wire [23:0] rounding_io_in_frac; // @[FPU.scala 274:24]
  wire  rounding_io_in_sign; // @[FPU.scala 274:24]
  wire  rounding_io_in_guard; // @[FPU.scala 274:24]
  wire  rounding_io_in_round; // @[FPU.scala 274:24]
  wire  rounding_io_in_sticky; // @[FPU.scala 274:24]
  wire [23:0] rounding_io_out_fracRounded; // @[FPU.scala 274:24]
  wire  rounding_io_out_fracCout; // @[FPU.scala 274:24]
  reg  REG; // @[util.scala 104:58]
  reg  REG_1; // @[util.scala 104:58]
  reg  REG_2; // @[util.scala 104:58]
  reg  REG_3; // @[util.scala 104:58]
  reg  REG_4; // @[util.scala 104:58]
  wire  _T_5 = ~io_out_ready & (REG & REG_1 & REG_2 & REG_3 & REG_4); // @[util.scala 106:26]
  wire  _T_6 = ~(~io_out_ready & (REG & REG_1 & REG_2 & REG_3 & REG_4)); // @[util.scala 106:10]
  wire  _T_12 = ~(~io_out_ready & (REG_1 & REG_2 & REG_3 & REG_4)); // @[util.scala 106:10]
  wire  _T_17 = ~(~io_out_ready & (REG_2 & REG_3 & REG_4)); // @[util.scala 106:10]
  wire  _T_21 = ~(~io_out_ready & (REG_3 & REG_4)); // @[util.scala 106:10]
  wire  _T_24 = ~(~io_out_ready & REG_4); // @[util.scala 106:10]
  wire [31:0] _a_x_T_2 = io_in_bits_op[1] ? 32'h0 : io_in_bits_b; // @[FPU.scala 87:10]
  wire [31:0] a_x = io_in_bits_op[2] ? io_in_bits_c : _a_x_T_2; // @[FPU.scala 85:16]
  wire  a_sign = a_x[31] ^ io_in_bits_op[0]; // @[FPU.scala 92:26]
  wire [31:0] a = {a_sign,a_x[30:0]}; // @[Cat.scala 31:58]
  wire [31:0] c = io_in_bits_op[2:1] == 2'h0 ? 32'h3f800000 : io_in_bits_b; // @[FPU.scala 96:14]
  wire [22:0] f32_frac = a[22:0]; // @[util.scala 46:46]
  wire [7:0] f32_exp = a[30:23]; // @[util.scala 46:46]
  wire  f32_sign = a[31]; // @[util.scala 46:46]
  wire [8:0] _exp_T_1 = {1'h0,f32_exp}; // @[util.scala 76:47]
  wire [8:0] _exp_T_7 = $signed(_exp_T_1) - 9'sh7f; // @[FPU.scala 106:22]
  wire [8:0] e = Classify_io_isSubnormal ? $signed(-9'sh7e) : $signed(_exp_T_7); // @[FPU.scala 104:18]
  wire  _fracExt_T = ~Classify_io_isSubnormal; // @[FPU.scala 108:40]
  wire [23:0] _fracExt_T_1 = {_fracExt_T,f32_frac}; // @[Cat.scala 31:58]
  wire [22:0] f32_1_frac = io_in_bits_a[22:0]; // @[util.scala 46:46]
  wire [7:0] f32_1_exp = io_in_bits_a[30:23]; // @[util.scala 46:46]
  wire  f32_1_sign = io_in_bits_a[31]; // @[util.scala 46:46]
  wire [8:0] _exp_T_9 = {1'h0,f32_1_exp}; // @[util.scala 76:47]
  wire [8:0] _exp_T_15 = $signed(_exp_T_9) - 9'sh7f; // @[FPU.scala 106:22]
  wire [8:0] e_1 = Classify_1_io_isSubnormal ? $signed(-9'sh7e) : $signed(_exp_T_15); // @[FPU.scala 104:18]
  wire  _fracExt_T_2 = ~Classify_1_io_isSubnormal; // @[FPU.scala 108:40]
  wire [23:0] _fracExt_T_3 = {_fracExt_T_2,f32_1_frac}; // @[Cat.scala 31:58]
  wire [23:0] f_1 = Classify_1_io_isZero ? 24'h0 : _fracExt_T_3; // @[FPU.scala 108:22]
  wire [22:0] f32_2_frac = c[22:0]; // @[util.scala 46:46]
  wire [7:0] f32_2_exp = c[30:23]; // @[util.scala 46:46]
  wire  f32_2_sign = c[31]; // @[util.scala 46:46]
  wire [8:0] _exp_T_17 = {1'h0,f32_2_exp}; // @[util.scala 76:47]
  wire [8:0] _exp_T_23 = $signed(_exp_T_17) - 9'sh7f; // @[FPU.scala 106:22]
  wire [8:0] e_2 = Classify_2_io_isSubnormal ? $signed(-9'sh7e) : $signed(_exp_T_23); // @[FPU.scala 104:18]
  wire  _fracExt_T_4 = ~Classify_2_io_isSubnormal; // @[FPU.scala 108:40]
  wire [23:0] _fracExt_T_5 = {_fracExt_T_4,f32_2_frac}; // @[Cat.scala 31:58]
  wire [23:0] f_2 = Classify_2_io_isZero ? 24'h0 : _fracExt_T_5; // @[FPU.scala 108:22]
  wire  prodIsZero = Classify_1_io_isZero | Classify_2_io_isZero; // @[FPU.scala 123:44]
  wire  prodSign = f32_1_sign ^ f32_2_sign ^ io_in_bits_op[2:1] == 2'h3; // @[FPU.scala 124:45]
  wire [9:0] _WIRE_4 = {{1{e_1[8]}},e_1}; // @[FPU.scala 113:35 118:17]
  wire [9:0] _WIRE_5 = {{1{e_2[8]}},e_2}; // @[FPU.scala 113:35 118:17]
  wire [9:0] _prodExpRaw_T_2 = $signed(_WIRE_4) + $signed(_WIRE_5); // @[FPU.scala 127:13]
  wire [9:0] prodExpRaw = prodIsZero ? $signed(-10'sh7f) : $signed(_prodExpRaw_T_2); // @[FPU.scala 125:28]
  wire  _zeroResultSign_T_6 = f32_sign & prodSign | (f32_sign | prodSign) & io_in_bits_rm == 3'h2; // @[FPU.scala 132:27]
  wire  hasNaN = Classify_io_isNaN | Classify_1_io_isNaN | Classify_2_io_isNaN; // @[FPU.scala 135:47]
  wire  hasInf = Classify_io_isInf | Classify_1_io_isInf | Classify_2_io_isInf; // @[FPU.scala 139:35]
  wire  prodHasInf = Classify_1_io_isInf | Classify_2_io_isInf; // @[FPU.scala 140:30]
  wire  addInfInvalid = Classify_io_isInf & prodHasInf & (f32_sign ^ prodSign) & ~(Classify_io_isInf ^ prodHasInf); // @[FPU.scala 142:73]
  wire  zeroMulInf = prodIsZero & prodHasInf; // @[FPU.scala 143:36]
  wire  infInvalid = addInfInvalid | zeroMulInf; // @[FPU.scala 144:39]
  wire  specialCase = hasNaN | hasInf; // @[FPU.scala 146:32]
  wire  _specialOutput_T = hasNaN | infInvalid; // @[FPU.scala 148:13]
  wire [31:0] _specialOutput_T_7 = {f32_sign,31'h7f800000}; // @[Cat.scala 31:58]
  wire [31:0] _specialOutput_T_11 = {prodSign,31'h7f800000}; // @[Cat.scala 31:58]
  wire [9:0] prodExpAdj = $signed(prodExpRaw) + 10'sh1b; // @[FPU.scala 152:31]
  wire [9:0] _WIRE_3 = {{1{e[8]}},e}; // @[FPU.scala 113:35 118:17]
  wire [9:0] expDiff = $signed(prodExpAdj) - $signed(_WIRE_3); // @[FPU.scala 153:28]
  wire  _s1_rm_T_7 = io_in_valid & _T_6; // @[util.scala 109:84]
  reg [2:0] s1_rm; // @[Reg.scala 16:16]
  reg  s1_zeroSign; // @[Reg.scala 16:16]
  reg  s1_specialCase; // @[Reg.scala 16:16]
  reg [31:0] s1_specialOutput; // @[Reg.scala 16:16]
  reg  s1_aSign; // @[Reg.scala 16:16]
  reg [9:0] s1_aExpRaw; // @[Reg.scala 16:16]
  reg [23:0] s1_aFrac; // @[Reg.scala 16:16]
  reg  s1_prodSign; // @[Reg.scala 16:16]
  reg [9:0] s1_prodExpAdj; // @[Reg.scala 16:16]
  reg [9:0] s1_expDiff; // @[Reg.scala 16:16]
  wire  _s1_discardProdFrac_T_2 = prodIsZero | expDiff[9]; // @[FPU.scala 169:45]
  reg  s1_discardProdFrac; // @[Reg.scala 16:16]
  wire  _s1_discardAFrac_T_1 = Classify_io_isZero | $signed(expDiff) > 10'sh4d; // @[FPU.scala 170:50]
  reg  s1_discardAFrac; // @[Reg.scala 16:16]
  reg [49:0] s1_mult_sum; // @[Reg.scala 16:16]
  wire [9:0] _alignedAFrac_T_1 = s1_discardProdFrac ? 10'h0 : s1_expDiff; // @[FPU.scala 178:39]
  wire [76:0] alignedAFrac_x_ext = {s1_aFrac,53'h0}; // @[Cat.scala 31:58]
  wire [6:0] alignedAFrac_realShiftAmt = _alignedAFrac_T_1 > 10'h4c ? 7'h4d : _alignedAFrac_T_1[6:0]; // @[util.scala 125:27]
  wire [6:0] _alignedAFrac_mask_T_2 = 7'h4d - alignedAFrac_realShiftAmt; // @[util.scala 129:48]
  wire [76:0] alignedAFrac_mask = 77'h1fffffffffffffffffff >> _alignedAFrac_mask_T_2; // @[util.scala 129:41]
  wire [76:0] alignedAFrac_x_shifted = alignedAFrac_x_ext >> alignedAFrac_realShiftAmt; // @[util.scala 131:24]
  wire [76:0] _alignedAFrac_T_3 = alignedAFrac_mask & alignedAFrac_x_ext; // @[util.scala 132:32]
  wire [76:0] _GEN_65 = {{76'd0}, |_alignedAFrac_T_3}; // @[util.scala 132:23]
  wire [76:0] _alignedAFrac_T_5 = alignedAFrac_x_shifted | _GEN_65; // @[util.scala 132:23]
  wire [77:0] alignedAFrac = {1'h0,_alignedAFrac_T_5}; // @[Cat.scala 31:58]
  wire [77:0] alignedAFracNeg = 78'h0 - alignedAFrac; // @[FPU.scala 180:25]
  wire  effSub = s1_prodSign ^ s1_aSign; // @[FPU.scala 181:28]
  wire [49:0] _mul_prod_T_2 = {{1'd0}, s1_mult_sum[48:0]}; // @[FPU.scala 182:40]
  wire [48:0] mul_prod = _mul_prod_T_2[48:0]; // @[FPU.scala 182:40]
  wire  _expPreNorm_T_1 = s1_discardAFrac | ~s1_discardProdFrac; // @[FPU.scala 184:40]
  wire  _s2_rm_T_6 = REG & _T_12; // @[util.scala 109:84]
  reg [2:0] s2_rm; // @[Reg.scala 16:16]
  reg  s2_zeroSign; // @[Reg.scala 16:16]
  reg  s2_specialCase; // @[Reg.scala 16:16]
  reg [31:0] s2_specialOutput; // @[Reg.scala 16:16]
  reg  s2_aSign; // @[Reg.scala 16:16]
  reg  s2_prodSign; // @[Reg.scala 16:16]
  reg [9:0] s2_expPreNorm; // @[Reg.scala 16:16]
  reg [48:0] s2_prod; // @[Reg.scala 16:16]
  reg [77:0] s2_aFracNeg; // @[Reg.scala 16:16]
  reg [77:0] s2_aFrac; // @[Reg.scala 16:16]
  reg  s2_effSub; // @[Reg.scala 16:16]
  wire [51:0] _prodMinusA_T = {s2_prod,3'h0}; // @[Cat.scala 31:58]
  wire [77:0] _GEN_66 = {{26'd0}, _prodMinusA_T}; // @[FPU.scala 200:43]
  wire [77:0] prodMinusA = _GEN_66 + s2_aFracNeg; // @[FPU.scala 200:43]
  wire  prodMinusA_Sign = prodMinusA[77]; // @[FPU.scala 201:40]
  wire [77:0] aMinusProd = 78'h0 - prodMinusA; // @[FPU.scala 202:20]
  wire [77:0] prodAddA = _GEN_66 + s2_aFrac; // @[FPU.scala 203:41]
  wire [77:0] _res_T = prodMinusA_Sign ? aMinusProd : prodMinusA; // @[FPU.scala 206:8]
  wire [77:0] res = s2_effSub ? _res_T : prodAddA; // @[FPU.scala 205:16]
  wire  _resSign_T = ~prodMinusA_Sign; // @[FPU.scala 215:7]
  wire  _resSign_T_1 = s2_aSign | _resSign_T; // @[FPU.scala 213:8]
  wire  _resSign_T_2 = s2_aSign & prodMinusA_Sign; // @[FPU.scala 217:8]
  wire [76:0] fracPreNorm = res[76:0]; // @[FPU.scala 222:29]
  wire [6:0] _normShift_T_78 = fracPreNorm[1] ? 7'h4b : 7'h4c; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_79 = fracPreNorm[2] ? 7'h4a : _normShift_T_78; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_80 = fracPreNorm[3] ? 7'h49 : _normShift_T_79; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_81 = fracPreNorm[4] ? 7'h48 : _normShift_T_80; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_82 = fracPreNorm[5] ? 7'h47 : _normShift_T_81; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_83 = fracPreNorm[6] ? 7'h46 : _normShift_T_82; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_84 = fracPreNorm[7] ? 7'h45 : _normShift_T_83; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_85 = fracPreNorm[8] ? 7'h44 : _normShift_T_84; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_86 = fracPreNorm[9] ? 7'h43 : _normShift_T_85; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_87 = fracPreNorm[10] ? 7'h42 : _normShift_T_86; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_88 = fracPreNorm[11] ? 7'h41 : _normShift_T_87; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_89 = fracPreNorm[12] ? 7'h40 : _normShift_T_88; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_90 = fracPreNorm[13] ? 7'h3f : _normShift_T_89; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_91 = fracPreNorm[14] ? 7'h3e : _normShift_T_90; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_92 = fracPreNorm[15] ? 7'h3d : _normShift_T_91; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_93 = fracPreNorm[16] ? 7'h3c : _normShift_T_92; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_94 = fracPreNorm[17] ? 7'h3b : _normShift_T_93; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_95 = fracPreNorm[18] ? 7'h3a : _normShift_T_94; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_96 = fracPreNorm[19] ? 7'h39 : _normShift_T_95; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_97 = fracPreNorm[20] ? 7'h38 : _normShift_T_96; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_98 = fracPreNorm[21] ? 7'h37 : _normShift_T_97; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_99 = fracPreNorm[22] ? 7'h36 : _normShift_T_98; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_100 = fracPreNorm[23] ? 7'h35 : _normShift_T_99; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_101 = fracPreNorm[24] ? 7'h34 : _normShift_T_100; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_102 = fracPreNorm[25] ? 7'h33 : _normShift_T_101; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_103 = fracPreNorm[26] ? 7'h32 : _normShift_T_102; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_104 = fracPreNorm[27] ? 7'h31 : _normShift_T_103; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_105 = fracPreNorm[28] ? 7'h30 : _normShift_T_104; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_106 = fracPreNorm[29] ? 7'h2f : _normShift_T_105; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_107 = fracPreNorm[30] ? 7'h2e : _normShift_T_106; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_108 = fracPreNorm[31] ? 7'h2d : _normShift_T_107; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_109 = fracPreNorm[32] ? 7'h2c : _normShift_T_108; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_110 = fracPreNorm[33] ? 7'h2b : _normShift_T_109; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_111 = fracPreNorm[34] ? 7'h2a : _normShift_T_110; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_112 = fracPreNorm[35] ? 7'h29 : _normShift_T_111; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_113 = fracPreNorm[36] ? 7'h28 : _normShift_T_112; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_114 = fracPreNorm[37] ? 7'h27 : _normShift_T_113; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_115 = fracPreNorm[38] ? 7'h26 : _normShift_T_114; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_116 = fracPreNorm[39] ? 7'h25 : _normShift_T_115; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_117 = fracPreNorm[40] ? 7'h24 : _normShift_T_116; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_118 = fracPreNorm[41] ? 7'h23 : _normShift_T_117; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_119 = fracPreNorm[42] ? 7'h22 : _normShift_T_118; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_120 = fracPreNorm[43] ? 7'h21 : _normShift_T_119; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_121 = fracPreNorm[44] ? 7'h20 : _normShift_T_120; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_122 = fracPreNorm[45] ? 7'h1f : _normShift_T_121; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_123 = fracPreNorm[46] ? 7'h1e : _normShift_T_122; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_124 = fracPreNorm[47] ? 7'h1d : _normShift_T_123; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_125 = fracPreNorm[48] ? 7'h1c : _normShift_T_124; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_126 = fracPreNorm[49] ? 7'h1b : _normShift_T_125; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_127 = fracPreNorm[50] ? 7'h1a : _normShift_T_126; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_128 = fracPreNorm[51] ? 7'h19 : _normShift_T_127; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_129 = fracPreNorm[52] ? 7'h18 : _normShift_T_128; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_130 = fracPreNorm[53] ? 7'h17 : _normShift_T_129; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_131 = fracPreNorm[54] ? 7'h16 : _normShift_T_130; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_132 = fracPreNorm[55] ? 7'h15 : _normShift_T_131; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_133 = fracPreNorm[56] ? 7'h14 : _normShift_T_132; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_134 = fracPreNorm[57] ? 7'h13 : _normShift_T_133; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_135 = fracPreNorm[58] ? 7'h12 : _normShift_T_134; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_136 = fracPreNorm[59] ? 7'h11 : _normShift_T_135; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_137 = fracPreNorm[60] ? 7'h10 : _normShift_T_136; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_138 = fracPreNorm[61] ? 7'hf : _normShift_T_137; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_139 = fracPreNorm[62] ? 7'he : _normShift_T_138; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_140 = fracPreNorm[63] ? 7'hd : _normShift_T_139; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_141 = fracPreNorm[64] ? 7'hc : _normShift_T_140; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_142 = fracPreNorm[65] ? 7'hb : _normShift_T_141; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_143 = fracPreNorm[66] ? 7'ha : _normShift_T_142; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_144 = fracPreNorm[67] ? 7'h9 : _normShift_T_143; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_145 = fracPreNorm[68] ? 7'h8 : _normShift_T_144; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_146 = fracPreNorm[69] ? 7'h7 : _normShift_T_145; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_147 = fracPreNorm[70] ? 7'h6 : _normShift_T_146; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_148 = fracPreNorm[71] ? 7'h5 : _normShift_T_147; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_149 = fracPreNorm[72] ? 7'h4 : _normShift_T_148; // @[Mux.scala 47:70]
  wire [6:0] _normShift_T_150 = fracPreNorm[73] ? 7'h3 : _normShift_T_149; // @[Mux.scala 47:70]
  wire  _s3_ovSetInf_T_5 = REG_1 & _T_17; // @[util.scala 109:84]
  reg [2:0] s3_rm; // @[Reg.scala 16:16]
  reg  s3_zeroSign; // @[Reg.scala 16:16]
  reg  s3_specialCase; // @[Reg.scala 16:16]
  reg [31:0] s3_specialOutput; // @[Reg.scala 16:16]
  reg  s3_resSign; // @[Reg.scala 16:16]
  reg [76:0] s3_fracPreNorm; // @[Reg.scala 16:16]
  reg [9:0] s3_expPreNorm; // @[Reg.scala 16:16]
  reg [6:0] s3_normShift; // @[Reg.scala 16:16]
  wire [7:0] _expPostNorm_T_1 = {1'h0,s3_normShift}; // @[util.scala 76:47]
  wire [9:0] _GEN_68 = {{2{_expPostNorm_T_1[7]}},_expPostNorm_T_1}; // @[FPU.scala 247:35]
  wire [9:0] expPostNorm = $signed(s3_expPreNorm) - $signed(_GEN_68); // @[FPU.scala 247:35]
  wire [9:0] denormShift = -10'sh7e - $signed(expPostNorm); // @[FPU.scala 248:47]
  wire [9:0] _leftShift_T_4 = denormShift[9] ? $signed(10'sh0) : $signed(denormShift); // @[FPU.scala 250:44]
  wire [9:0] rightShift = $signed(denormShift) - $signed(_GEN_68); // @[FPU.scala 251:32]
  wire [9:0] _fracShifted_T_2 = $signed(_GEN_68) - $signed(_leftShift_T_4); // @[FPU.scala 253:50]
  wire [203:0] _GEN_5 = {{127'd0}, s3_fracPreNorm}; // @[util.scala 141:9]
  wire [203:0] _fracShifted_x_shifted_T_2 = _GEN_5 << _fracShifted_T_2[6:0]; // @[util.scala 141:9]
  wire [203:0] _fracShifted_x_shifted_T_3 = _fracShifted_T_2 > 10'h4c ? 204'h0 : _fracShifted_x_shifted_T_2; // @[util.scala 139:21]
  wire [76:0] fracShifted_x_shifted = _fracShifted_x_shifted_T_3[76:0]; // @[util.scala 138:25 139:15]
  wire [26:0] _GEN_71 = {{26'd0}, |fracShifted_x_shifted[49:0]}; // @[util.scala 143:23]
  wire [26:0] _fracShifted_T_6 = fracShifted_x_shifted[76:50] | _GEN_71; // @[util.scala 143:23]
  wire [9:0] _fracShifted_T_7 = $signed(denormShift) - $signed(_GEN_68); // @[FPU.scala 254:52]
  wire [4:0] fracShifted_realShiftAmt = _fracShifted_T_7 > 10'h1a ? 5'h1b : _fracShifted_T_7[4:0]; // @[util.scala 125:27]
  wire [4:0] _fracShifted_mask_T_2 = 5'h1b - fracShifted_realShiftAmt; // @[util.scala 129:48]
  wire [76:0] fracShifted_mask = 77'h1fffffffffffffffffff >> _fracShifted_mask_T_2; // @[util.scala 129:41]
  wire [76:0] fracShifted_x_shifted_1 = s3_fracPreNorm >> fracShifted_realShiftAmt; // @[util.scala 131:24]
  wire [76:0] _fracShifted_T_9 = fracShifted_mask & s3_fracPreNorm; // @[util.scala 132:32]
  wire [26:0] _GEN_72 = {{26'd0}, |_fracShifted_T_9}; // @[util.scala 132:23]
  wire [26:0] _fracShifted_T_11 = fracShifted_x_shifted_1[76:50] | _GEN_72; // @[util.scala 132:23]
  wire  _s4_rm_T_4 = REG_2 & _T_21; // @[util.scala 109:84]
  reg [2:0] s4_rm; // @[Reg.scala 16:16]
  reg  s4_zeroSign; // @[Reg.scala 16:16]
  reg  s4_specialCase; // @[Reg.scala 16:16]
  reg [31:0] s4_specialOutput; // @[Reg.scala 16:16]
  reg  s4_resSign; // @[Reg.scala 16:16]
  reg [26:0] s4_fracShifted; // @[Reg.scala 16:16]
  reg [9:0] s4_expPostNorm; // @[Reg.scala 16:16]
  reg [9:0] s4_denormShift; // @[Reg.scala 16:16]
  wire [23:0] fracUnrounded = s4_fracShifted[26:3]; // @[FPU.scala 270:42]
  wire  fracCout = ~fracUnrounded[23] ? rounding_io_out_fracRounded[23] : rounding_io_out_fracCout; // @[FPU.scala 283:21]
  wire [24:0] _isZeroResult_T = {fracCout,rounding_io_out_fracRounded}; // @[Cat.scala 31:58]
  wire  isZeroResult = ~(|_isZeroResult_T); // @[FPU.scala 288:22]
  wire [9:0] _expRounded_T_7 = $signed(s4_expPostNorm) + 10'sh7f; // @[FPU.scala 291:20]
  wire [9:0] _expRounded_T_8 = $signed(s4_denormShift) > 10'sh0 | isZeroResult ? $signed(10'sh0) : $signed(
    _expRounded_T_7); // @[FPU.scala 289:23]
  wire [1:0] _expRounded_T_10 = {1'h0,fracCout}; // @[util.scala 76:47]
  wire [9:0] _GEN_73 = {{8{_expRounded_T_10[1]}},_expRounded_T_10}; // @[FPU.scala 292:5]
  wire [9:0] expRounded = $signed(_expRounded_T_8) + $signed(_GEN_73); // @[FPU.scala 292:5]
  wire  _s5_sign_T_4 = REG_3 & _T_24; // @[util.scala 109:84]
  reg  s5_sign; // @[Reg.scala 16:16]
  reg [9:0] s5_exp; // @[Reg.scala 16:16]
  reg [23:0] s5_frac; // @[Reg.scala 16:16]
  reg  s5_specialCase; // @[Reg.scala 16:16]
  reg [31:0] s5_specialOutput; // @[Reg.scala 16:16]
  wire [31:0] commonResult = {s5_sign,s5_exp[7:0],s5_frac[22:0]}; // @[Cat.scala 31:58]
  Classify Classify ( // @[FPU.scala 99:38]
    .io_in(Classify_io_in),
    .io_isNegInf(Classify_io_isNegInf),
    .io_isNegNormal(Classify_io_isNegNormal),
    .io_isNegSubnormal(Classify_io_isNegSubnormal),
    .io_isNegZero(Classify_io_isNegZero),
    .io_isPosZero(Classify_io_isPosZero),
    .io_isPosSubnormal(Classify_io_isPosSubnormal),
    .io_isPosNormal(Classify_io_isPosNormal),
    .io_isPosInf(Classify_io_isPosInf),
    .io_isSNaN(Classify_io_isSNaN),
    .io_isQNaN(Classify_io_isQNaN),
    .io_isNaN(Classify_io_isNaN),
    .io_isInf(Classify_io_isInf),
    .io_isInfOrNaN(Classify_io_isInfOrNaN),
    .io_isSubnormal(Classify_io_isSubnormal),
    .io_isZero(Classify_io_isZero),
    .io_isSubnormalOrZero(Classify_io_isSubnormalOrZero)
  );
  Classify Classify_1 ( // @[FPU.scala 99:38]
    .io_in(Classify_1_io_in),
    .io_isNegInf(Classify_1_io_isNegInf),
    .io_isNegNormal(Classify_1_io_isNegNormal),
    .io_isNegSubnormal(Classify_1_io_isNegSubnormal),
    .io_isNegZero(Classify_1_io_isNegZero),
    .io_isPosZero(Classify_1_io_isPosZero),
    .io_isPosSubnormal(Classify_1_io_isPosSubnormal),
    .io_isPosNormal(Classify_1_io_isPosNormal),
    .io_isPosInf(Classify_1_io_isPosInf),
    .io_isSNaN(Classify_1_io_isSNaN),
    .io_isQNaN(Classify_1_io_isQNaN),
    .io_isNaN(Classify_1_io_isNaN),
    .io_isInf(Classify_1_io_isInf),
    .io_isInfOrNaN(Classify_1_io_isInfOrNaN),
    .io_isSubnormal(Classify_1_io_isSubnormal),
    .io_isZero(Classify_1_io_isZero),
    .io_isSubnormalOrZero(Classify_1_io_isSubnormalOrZero)
  );
  Classify Classify_2 ( // @[FPU.scala 99:38]
    .io_in(Classify_2_io_in),
    .io_isNegInf(Classify_2_io_isNegInf),
    .io_isNegNormal(Classify_2_io_isNegNormal),
    .io_isNegSubnormal(Classify_2_io_isNegSubnormal),
    .io_isNegZero(Classify_2_io_isNegZero),
    .io_isPosZero(Classify_2_io_isPosZero),
    .io_isPosSubnormal(Classify_2_io_isPosSubnormal),
    .io_isPosNormal(Classify_2_io_isPosNormal),
    .io_isPosInf(Classify_2_io_isPosInf),
    .io_isSNaN(Classify_2_io_isSNaN),
    .io_isQNaN(Classify_2_io_isQNaN),
    .io_isNaN(Classify_2_io_isNaN),
    .io_isInf(Classify_2_io_isInf),
    .io_isInfOrNaN(Classify_2_io_isInfOrNaN),
    .io_isSubnormal(Classify_2_io_isSubnormal),
    .io_isZero(Classify_2_io_isZero),
    .io_isSubnormalOrZero(Classify_2_io_isSubnormalOrZero)
  );
  ArrayMultiplier mult ( // @[FPU.scala 155:20]
    .io_a(mult_io_a),
    .io_b(mult_io_b),
    .io_sum(mult_io_sum)
  );
  RoundingUnit rounding ( // @[FPU.scala 274:24]
    .io_in_rm(rounding_io_in_rm),
    .io_in_frac(rounding_io_in_frac),
    .io_in_sign(rounding_io_in_sign),
    .io_in_guard(rounding_io_in_guard),
    .io_in_round(rounding_io_in_round),
    .io_in_sticky(rounding_io_in_sticky),
    .io_out_fracRounded(rounding_io_out_fracRounded),
    .io_out_fracCout(rounding_io_out_fracCout)
  );
  assign io_in_ready = ~_T_5; // @[util.scala 116:18]
  assign io_out_valid = REG_4; // @[util.scala 117:16]
  assign io_out_bits_result = s5_specialCase ? s5_specialOutput : commonResult; // @[FPU.scala 320:19]
  assign Classify_io_in = {a_sign,a_x[30:0]}; // @[Cat.scala 31:58]
  assign Classify_1_io_in = io_in_bits_a; // @[FPU.scala 100:60]
  assign Classify_2_io_in = io_in_bits_op[2:1] == 2'h0 ? 32'h3f800000 : io_in_bits_b; // @[FPU.scala 96:14]
  assign mult_io_a = {{1'd0}, f_1}; // @[FPU.scala 156:13]
  assign mult_io_b = {{1'd0}, f_2}; // @[FPU.scala 157:13]
  assign rounding_io_in_rm = s4_rm; // @[FPU.scala 275:21]
  assign rounding_io_in_frac = s4_fracShifted[26:3]; // @[FPU.scala 270:42]
  assign rounding_io_in_sign = s4_resSign; // @[FPU.scala 277:23]
  assign rounding_io_in_guard = s4_fracShifted[2]; // @[FPU.scala 271:49]
  assign rounding_io_in_round = s4_fracShifted[1]; // @[FPU.scala 272:51]
  assign rounding_io_in_sticky = |s4_fracShifted[0]; // @[FPU.scala 273:50]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 104:58]
      REG <= 1'h0; // @[util.scala 104:58]
    end else if (~(~io_out_ready & (REG & REG_1 & REG_2 & REG_3 & REG_4))) begin // @[util.scala 106:59]
      REG <= io_in_valid; // @[util.scala 106:71]
    end
    if (reset) begin // @[util.scala 104:58]
      REG_1 <= 1'h0; // @[util.scala 104:58]
    end else if (~(~io_out_ready & (REG_1 & REG_2 & REG_3 & REG_4))) begin // @[util.scala 106:59]
      REG_1 <= REG; // @[util.scala 106:71]
    end
    if (reset) begin // @[util.scala 104:58]
      REG_2 <= 1'h0; // @[util.scala 104:58]
    end else if (~(~io_out_ready & (REG_2 & REG_3 & REG_4))) begin // @[util.scala 106:59]
      REG_2 <= REG_1; // @[util.scala 106:71]
    end
    if (reset) begin // @[util.scala 104:58]
      REG_3 <= 1'h0; // @[util.scala 104:58]
    end else if (~(~io_out_ready & (REG_3 & REG_4))) begin // @[util.scala 106:59]
      REG_3 <= REG_2; // @[util.scala 106:71]
    end
    if (reset) begin // @[util.scala 104:58]
      REG_4 <= 1'h0; // @[util.scala 104:58]
    end else if (~(~io_out_ready & REG_4)) begin // @[util.scala 106:59]
      REG_4 <= REG_3; // @[util.scala 106:71]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_rm <= io_in_bits_rm; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      if (io_in_bits_op[2:1] == 2'h1) begin // @[FPU.scala 130:27]
        s1_zeroSign <= prodSign;
      end else begin
        s1_zeroSign <= _zeroResultSign_T_6;
      end
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_specialCase <= specialCase; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      if (_specialOutput_T) begin // @[Mux.scala 47:70]
        s1_specialOutput <= 32'h7fc00000;
      end else if (Classify_io_isInf) begin // @[Mux.scala 47:70]
        s1_specialOutput <= _specialOutput_T_7;
      end else begin
        s1_specialOutput <= _specialOutput_T_11;
      end
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_aSign <= f32_sign; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_aExpRaw <= _WIRE_3; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      if (Classify_io_isZero) begin // @[FPU.scala 108:22]
        s1_aFrac <= 24'h0;
      end else begin
        s1_aFrac <= _fracExt_T_1;
      end
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_prodSign <= prodSign; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_prodExpAdj <= prodExpAdj; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_expDiff <= expDiff; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_discardProdFrac <= _s1_discardProdFrac_T_2; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_discardAFrac <= _s1_discardAFrac_T_1; // @[Reg.scala 17:22]
    end
    if (_s1_rm_T_7) begin // @[Reg.scala 17:18]
      s1_mult_sum <= mult_io_sum; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_rm <= s1_rm; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_zeroSign <= s1_zeroSign; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_specialCase <= s1_specialCase; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_specialOutput <= s1_specialOutput; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_aSign <= s1_aSign; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_prodSign <= s1_prodSign; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      if (_expPreNorm_T_1) begin // @[FPU.scala 192:32]
        s2_expPreNorm <= s1_prodExpAdj;
      end else begin
        s2_expPreNorm <= s1_aExpRaw;
      end
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_prod <= mul_prod; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_aFracNeg <= alignedAFracNeg; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_aFrac <= alignedAFrac; // @[Reg.scala 17:22]
    end
    if (_s2_rm_T_6) begin // @[Reg.scala 17:18]
      s2_effSub <= effSub; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      s3_rm <= s2_rm; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      s3_zeroSign <= s2_zeroSign; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      s3_specialCase <= s2_specialCase; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      s3_specialOutput <= s2_specialOutput; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      if (s2_prodSign) begin // @[FPU.scala 212:20]
        s3_resSign <= _resSign_T_1;
      end else begin
        s3_resSign <= _resSign_T_2;
      end
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      s3_fracPreNorm <= fracPreNorm; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      s3_expPreNorm <= s2_expPreNorm; // @[Reg.scala 17:22]
    end
    if (_s3_ovSetInf_T_5) begin // @[Reg.scala 17:18]
      if (fracPreNorm[76]) begin // @[Mux.scala 47:70]
        s3_normShift <= 7'h0;
      end else if (fracPreNorm[75]) begin // @[Mux.scala 47:70]
        s3_normShift <= 7'h1;
      end else if (fracPreNorm[74]) begin // @[Mux.scala 47:70]
        s3_normShift <= 7'h2;
      end else begin
        s3_normShift <= _normShift_T_150;
      end
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_rm <= s3_rm; // @[Reg.scala 17:22]
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_zeroSign <= s3_zeroSign; // @[Reg.scala 17:22]
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_specialCase <= s3_specialCase; // @[Reg.scala 17:22]
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_specialOutput <= s3_specialOutput; // @[Reg.scala 17:22]
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_resSign <= s3_resSign; // @[Reg.scala 17:22]
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      if (rightShift[9]) begin // @[FPU.scala 252:24]
        s4_fracShifted <= _fracShifted_T_6;
      end else begin
        s4_fracShifted <= _fracShifted_T_11;
      end
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_expPostNorm <= expPostNorm; // @[Reg.scala 17:22]
    end
    if (_s4_rm_T_4) begin // @[Reg.scala 17:18]
      s4_denormShift <= denormShift; // @[Reg.scala 17:22]
    end
    if (_s5_sign_T_4) begin // @[Reg.scala 17:18]
      if (isZeroResult) begin // @[FPU.scala 304:26]
        s5_sign <= s4_zeroSign;
      end else begin
        s5_sign <= s4_resSign;
      end
    end
    if (_s5_sign_T_4) begin // @[Reg.scala 17:18]
      s5_exp <= expRounded; // @[Reg.scala 17:22]
    end
    if (_s5_sign_T_4) begin // @[Reg.scala 17:18]
      s5_frac <= rounding_io_out_fracRounded; // @[Reg.scala 17:22]
    end
    if (_s5_sign_T_4) begin // @[Reg.scala 17:18]
      s5_specialCase <= s4_specialCase; // @[Reg.scala 17:22]
    end
    if (_s5_sign_T_4) begin // @[Reg.scala 17:18]
      s5_specialOutput <= s4_specialOutput; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s1_rm = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  s1_zeroSign = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s1_specialCase = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s1_specialOutput = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  s1_aSign = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  s1_aExpRaw = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  s1_aFrac = _RAND_11[23:0];
  _RAND_12 = {1{`RANDOM}};
  s1_prodSign = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  s1_prodExpAdj = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  s1_expDiff = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  s1_discardProdFrac = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  s1_discardAFrac = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  s1_mult_sum = _RAND_17[49:0];
  _RAND_18 = {1{`RANDOM}};
  s2_rm = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  s2_zeroSign = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  s2_specialCase = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s2_specialOutput = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  s2_aSign = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  s2_prodSign = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  s2_expPreNorm = _RAND_24[9:0];
  _RAND_25 = {2{`RANDOM}};
  s2_prod = _RAND_25[48:0];
  _RAND_26 = {3{`RANDOM}};
  s2_aFracNeg = _RAND_26[77:0];
  _RAND_27 = {3{`RANDOM}};
  s2_aFrac = _RAND_27[77:0];
  _RAND_28 = {1{`RANDOM}};
  s2_effSub = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  s3_rm = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  s3_zeroSign = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  s3_specialCase = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  s3_specialOutput = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  s3_resSign = _RAND_33[0:0];
  _RAND_34 = {3{`RANDOM}};
  s3_fracPreNorm = _RAND_34[76:0];
  _RAND_35 = {1{`RANDOM}};
  s3_expPreNorm = _RAND_35[9:0];
  _RAND_36 = {1{`RANDOM}};
  s3_normShift = _RAND_36[6:0];
  _RAND_37 = {1{`RANDOM}};
  s4_rm = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  s4_zeroSign = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  s4_specialCase = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  s4_specialOutput = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  s4_resSign = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  s4_fracShifted = _RAND_42[26:0];
  _RAND_43 = {1{`RANDOM}};
  s4_expPostNorm = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  s4_denormShift = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  s5_sign = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  s5_exp = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  s5_frac = _RAND_47[23:0];
  _RAND_48 = {1{`RANDOM}};
  s5_specialCase = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  s5_specialOutput = _RAND_49[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_result,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_result
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_result [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_result_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_result_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_result_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_result_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_result_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_result_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_result_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_result_io_deq_bits_MPORT_en = 1'h1;
  assign ram_result_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_result_io_deq_bits_MPORT_data = ram_result[ram_result_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_result_MPORT_data = io_enq_bits_result;
  assign ram_result_MPORT_addr = 1'h0;
  assign ram_result_MPORT_mask = 1'h1;
  assign ram_result_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_result = ram_result_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_result_MPORT_en & ram_result_MPORT_mask) begin
      ram_result[ram_result_MPORT_addr] <= ram_result_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_result[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPU_CMP(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_op,
  input  [31:0] io_in_bits_a,
  input  [31:0] io_in_bits_b,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result
);
  wire [31:0] Classify_io_in; // @[FPU.scala 353:38]
  wire  Classify_io_isNegInf; // @[FPU.scala 353:38]
  wire  Classify_io_isNegNormal; // @[FPU.scala 353:38]
  wire  Classify_io_isNegSubnormal; // @[FPU.scala 353:38]
  wire  Classify_io_isNegZero; // @[FPU.scala 353:38]
  wire  Classify_io_isPosZero; // @[FPU.scala 353:38]
  wire  Classify_io_isPosSubnormal; // @[FPU.scala 353:38]
  wire  Classify_io_isPosNormal; // @[FPU.scala 353:38]
  wire  Classify_io_isPosInf; // @[FPU.scala 353:38]
  wire  Classify_io_isSNaN; // @[FPU.scala 353:38]
  wire  Classify_io_isQNaN; // @[FPU.scala 353:38]
  wire  Classify_io_isNaN; // @[FPU.scala 353:38]
  wire  Classify_io_isInf; // @[FPU.scala 353:38]
  wire  Classify_io_isInfOrNaN; // @[FPU.scala 353:38]
  wire  Classify_io_isSubnormal; // @[FPU.scala 353:38]
  wire  Classify_io_isZero; // @[FPU.scala 353:38]
  wire  Classify_io_isSubnormalOrZero; // @[FPU.scala 353:38]
  wire [31:0] Classify_1_io_in; // @[FPU.scala 353:38]
  wire  Classify_1_io_isNegInf; // @[FPU.scala 353:38]
  wire  Classify_1_io_isNegNormal; // @[FPU.scala 353:38]
  wire  Classify_1_io_isNegSubnormal; // @[FPU.scala 353:38]
  wire  Classify_1_io_isNegZero; // @[FPU.scala 353:38]
  wire  Classify_1_io_isPosZero; // @[FPU.scala 353:38]
  wire  Classify_1_io_isPosSubnormal; // @[FPU.scala 353:38]
  wire  Classify_1_io_isPosNormal; // @[FPU.scala 353:38]
  wire  Classify_1_io_isPosInf; // @[FPU.scala 353:38]
  wire  Classify_1_io_isSNaN; // @[FPU.scala 353:38]
  wire  Classify_1_io_isQNaN; // @[FPU.scala 353:38]
  wire  Classify_1_io_isNaN; // @[FPU.scala 353:38]
  wire  Classify_1_io_isInf; // @[FPU.scala 353:38]
  wire  Classify_1_io_isInfOrNaN; // @[FPU.scala 353:38]
  wire  Classify_1_io_isSubnormal; // @[FPU.scala 353:38]
  wire  Classify_1_io_isZero; // @[FPU.scala 353:38]
  wire  Classify_1_io_isSubnormalOrZero; // @[FPU.scala 353:38]
  wire  result_clock; // @[FPU.scala 395:20]
  wire  result_reset; // @[FPU.scala 395:20]
  wire  result_io_enq_ready; // @[FPU.scala 395:20]
  wire  result_io_enq_valid; // @[FPU.scala 395:20]
  wire [31:0] result_io_enq_bits_result; // @[FPU.scala 395:20]
  wire  result_io_deq_ready; // @[FPU.scala 395:20]
  wire  result_io_deq_valid; // @[FPU.scala 395:20]
  wire [31:0] result_io_deq_bits_result; // @[FPU.scala 395:20]
  wire  sign_0 = io_in_bits_a[31]; // @[FPU.scala 351:23]
  wire  sign_1 = io_in_bits_b[31]; // @[FPU.scala 351:23]
  wire [32:0] _subRes_T_1 = {1'h0,io_in_bits_a}; // @[util.scala 76:47]
  wire [32:0] _subRes_T_3 = {1'h0,io_in_bits_b}; // @[util.scala 76:47]
  wire [32:0] subRes = $signed(_subRes_T_1) - $signed(_subRes_T_3); // @[FPU.scala 352:30]
  wire  hasNaN = Classify_io_isNaN | Classify_1_io_isNaN; // @[FPU.scala 359:28]
  wire  bothNaN = Classify_io_isNaN & Classify_1_io_isNaN; // @[FPU.scala 360:29]
  wire  bothZero = io_in_bits_a[30:0] == 31'h0 & io_in_bits_b[30:0] == 31'h0; // @[FPU.scala 361:39]
  wire  uintEq = $signed(subRes) == 33'sh0; // @[FPU.scala 362:22]
  wire  uintLess = sign_0 ^ $signed(subRes) < 33'sh0; // @[FPU.scala 363:26]
  wire  eq = uintEq | bothZero; // @[FPU.scala 368:16]
  wire  _le_T = sign_0 != sign_1; // @[FPU.scala 369:20]
  wire  _le_T_1 = sign_0 | bothZero; // @[FPU.scala 370:13]
  wire  _le_T_2 = uintEq | uintLess; // @[FPU.scala 371:12]
  wire  le = sign_0 != sign_1 ? _le_T_1 : _le_T_2; // @[FPU.scala 369:12]
  wire  _lt_T_2 = sign_0 & ~bothZero; // @[FPU.scala 374:13]
  wire  _lt_T_4 = ~uintEq & uintLess; // @[FPU.scala 375:13]
  wire  lt = _le_T ? _lt_T_2 : _lt_T_4; // @[FPU.scala 373:12]
  wire  _fcmpResult_T_6 = io_in_bits_op[0] ? lt : le; // @[FPU.scala 379:58]
  wire  _fcmpResult_T_7 = io_in_bits_op[2] ? eq : _fcmpResult_T_6; // @[FPU.scala 379:43]
  wire  _fcmpResult_T_8 = io_in_bits_op[2] & io_in_bits_op[0] ? ~eq : _fcmpResult_T_7; // @[FPU.scala 379:23]
  wire [31:0] _fcmpResult_T_9 = {31'h0,_fcmpResult_T_8}; // @[Cat.scala 31:58]
  wire [31:0] fcmpResult = hasNaN ? 32'h0 : _fcmpResult_T_9; // @[FPU.scala 377:23]
  wire  _min_T_4 = lt | eq & sign_0; // @[FPU.scala 383:14]
  wire  _min_T_5 = ~Classify_io_isNaN; // @[FPU.scala 383:37]
  wire [31:0] _min_T_7 = (lt | eq & sign_0) & ~Classify_io_isNaN ? io_in_bits_a : io_in_bits_b; // @[FPU.scala 383:8]
  wire [31:0] min = bothNaN ? 32'h7fc00000 : _min_T_7; // @[FPU.scala 381:16]
  wire [31:0] _max_T_8 = ~_min_T_4 & _min_T_5 ? io_in_bits_a : io_in_bits_b; // @[FPU.scala 390:8]
  wire [31:0] max = bothNaN ? 32'h7fc00000 : _max_T_8; // @[FPU.scala 388:16]
  wire [31:0] _result_io_enq_bits_result_T_2 = io_in_bits_op == 3'h1 ? max : fcmpResult; // @[FPU.scala 396:54]
  Classify Classify ( // @[FPU.scala 353:38]
    .io_in(Classify_io_in),
    .io_isNegInf(Classify_io_isNegInf),
    .io_isNegNormal(Classify_io_isNegNormal),
    .io_isNegSubnormal(Classify_io_isNegSubnormal),
    .io_isNegZero(Classify_io_isNegZero),
    .io_isPosZero(Classify_io_isPosZero),
    .io_isPosSubnormal(Classify_io_isPosSubnormal),
    .io_isPosNormal(Classify_io_isPosNormal),
    .io_isPosInf(Classify_io_isPosInf),
    .io_isSNaN(Classify_io_isSNaN),
    .io_isQNaN(Classify_io_isQNaN),
    .io_isNaN(Classify_io_isNaN),
    .io_isInf(Classify_io_isInf),
    .io_isInfOrNaN(Classify_io_isInfOrNaN),
    .io_isSubnormal(Classify_io_isSubnormal),
    .io_isZero(Classify_io_isZero),
    .io_isSubnormalOrZero(Classify_io_isSubnormalOrZero)
  );
  Classify Classify_1 ( // @[FPU.scala 353:38]
    .io_in(Classify_1_io_in),
    .io_isNegInf(Classify_1_io_isNegInf),
    .io_isNegNormal(Classify_1_io_isNegNormal),
    .io_isNegSubnormal(Classify_1_io_isNegSubnormal),
    .io_isNegZero(Classify_1_io_isNegZero),
    .io_isPosZero(Classify_1_io_isPosZero),
    .io_isPosSubnormal(Classify_1_io_isPosSubnormal),
    .io_isPosNormal(Classify_1_io_isPosNormal),
    .io_isPosInf(Classify_1_io_isPosInf),
    .io_isSNaN(Classify_1_io_isSNaN),
    .io_isQNaN(Classify_1_io_isQNaN),
    .io_isNaN(Classify_1_io_isNaN),
    .io_isInf(Classify_1_io_isInf),
    .io_isInfOrNaN(Classify_1_io_isInfOrNaN),
    .io_isSubnormal(Classify_1_io_isSubnormal),
    .io_isZero(Classify_1_io_isZero),
    .io_isSubnormalOrZero(Classify_1_io_isSubnormalOrZero)
  );
  Queue_5 result ( // @[FPU.scala 395:20]
    .clock(result_clock),
    .reset(result_reset),
    .io_enq_ready(result_io_enq_ready),
    .io_enq_valid(result_io_enq_valid),
    .io_enq_bits_result(result_io_enq_bits_result),
    .io_deq_ready(result_io_deq_ready),
    .io_deq_valid(result_io_deq_valid),
    .io_deq_bits_result(result_io_deq_bits_result)
  );
  assign io_in_ready = result_io_enq_ready; // @[FPU.scala 403:14]
  assign io_out_valid = result_io_deq_valid; // @[FPU.scala 405:16]
  assign io_out_bits_result = result_io_deq_bits_result; // @[FPU.scala 406:14]
  assign Classify_io_in = io_in_bits_a; // @[FPU.scala 354:50]
  assign Classify_1_io_in = io_in_bits_b; // @[FPU.scala 354:50]
  assign result_clock = clock;
  assign result_reset = reset;
  assign result_io_enq_valid = io_in_valid; // @[FPU.scala 402:22]
  assign result_io_enq_bits_result = io_in_bits_op == 3'h0 ? min : _result_io_enq_bits_result_T_2; // @[FPU.scala 396:35]
  assign result_io_deq_ready = io_out_ready; // @[FPU.scala 407:22]
endmodule
module FPU_FMV(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_op,
  input  [31:0] io_in_bits_a,
  input  [31:0] io_in_bits_b,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result
);
  wire [31:0] Classify_io_in; // @[FPU.scala 541:19]
  wire  Classify_io_isNegInf; // @[FPU.scala 541:19]
  wire  Classify_io_isNegNormal; // @[FPU.scala 541:19]
  wire  Classify_io_isNegSubnormal; // @[FPU.scala 541:19]
  wire  Classify_io_isNegZero; // @[FPU.scala 541:19]
  wire  Classify_io_isPosZero; // @[FPU.scala 541:19]
  wire  Classify_io_isPosSubnormal; // @[FPU.scala 541:19]
  wire  Classify_io_isPosNormal; // @[FPU.scala 541:19]
  wire  Classify_io_isPosInf; // @[FPU.scala 541:19]
  wire  Classify_io_isSNaN; // @[FPU.scala 541:19]
  wire  Classify_io_isQNaN; // @[FPU.scala 541:19]
  wire  Classify_io_isNaN; // @[FPU.scala 541:19]
  wire  Classify_io_isInf; // @[FPU.scala 541:19]
  wire  Classify_io_isInfOrNaN; // @[FPU.scala 541:19]
  wire  Classify_io_isSubnormal; // @[FPU.scala 541:19]
  wire  Classify_io_isZero; // @[FPU.scala 541:19]
  wire  Classify_io_isSubnormalOrZero; // @[FPU.scala 541:19]
  wire  result_reg_clock; // @[FPU.scala 560:24]
  wire  result_reg_reset; // @[FPU.scala 560:24]
  wire  result_reg_io_enq_ready; // @[FPU.scala 560:24]
  wire  result_reg_io_enq_valid; // @[FPU.scala 560:24]
  wire [31:0] result_reg_io_enq_bits_result; // @[FPU.scala 560:24]
  wire  result_reg_io_deq_ready; // @[FPU.scala 560:24]
  wire  result_reg_io_deq_valid; // @[FPU.scala 560:24]
  wire [31:0] result_reg_io_deq_bits_result; // @[FPU.scala 560:24]
  wire  _sgnjSign_T_8 = io_in_bits_op[0] ? ~io_in_bits_b[31] : io_in_bits_a[31] ^ io_in_bits_b[31]; // @[FPU.scala 538:8]
  wire  sgnjSign = io_in_bits_op[1] ? io_in_bits_b[31] : _sgnjSign_T_8; // @[FPU.scala 536:21]
  wire  resSign = io_in_bits_op[2] ? sgnjSign : io_in_bits_a[31]; // @[FPU.scala 540:20]
  wire [9:0] classifyResult = {Classify_io_isQNaN,Classify_io_isSNaN,Classify_io_isPosInf,Classify_io_isPosNormal,
    Classify_io_isPosSubnormal,Classify_io_isPosZero,Classify_io_isNegZero,Classify_io_isNegSubnormal,
    Classify_io_isNegNormal,Classify_io_isNegInf}; // @[Cat.scala 31:58]
  wire [31:0] _result_T_2 = {resSign,io_in_bits_a[30:0]}; // @[Cat.scala 31:58]
  Classify Classify ( // @[FPU.scala 541:19]
    .io_in(Classify_io_in),
    .io_isNegInf(Classify_io_isNegInf),
    .io_isNegNormal(Classify_io_isNegNormal),
    .io_isNegSubnormal(Classify_io_isNegSubnormal),
    .io_isNegZero(Classify_io_isNegZero),
    .io_isPosZero(Classify_io_isPosZero),
    .io_isPosSubnormal(Classify_io_isPosSubnormal),
    .io_isPosNormal(Classify_io_isPosNormal),
    .io_isPosInf(Classify_io_isPosInf),
    .io_isSNaN(Classify_io_isSNaN),
    .io_isQNaN(Classify_io_isQNaN),
    .io_isNaN(Classify_io_isNaN),
    .io_isInf(Classify_io_isInf),
    .io_isInfOrNaN(Classify_io_isInfOrNaN),
    .io_isSubnormal(Classify_io_isSubnormal),
    .io_isZero(Classify_io_isZero),
    .io_isSubnormalOrZero(Classify_io_isSubnormalOrZero)
  );
  Queue_5 result_reg ( // @[FPU.scala 560:24]
    .clock(result_reg_clock),
    .reset(result_reg_reset),
    .io_enq_ready(result_reg_io_enq_ready),
    .io_enq_valid(result_reg_io_enq_valid),
    .io_enq_bits_result(result_reg_io_enq_bits_result),
    .io_deq_ready(result_reg_io_deq_ready),
    .io_deq_valid(result_reg_io_deq_valid),
    .io_deq_bits_result(result_reg_io_deq_bits_result)
  );
  assign io_in_ready = result_reg_io_enq_ready; // @[FPU.scala 564:14]
  assign io_out_valid = result_reg_io_deq_valid; // @[FPU.scala 566:16]
  assign io_out_bits_result = result_reg_io_deq_bits_result; // @[FPU.scala 567:14]
  assign Classify_io_in = io_in_bits_a; // @[FPU.scala 542:10]
  assign result_reg_clock = clock;
  assign result_reg_reset = reset;
  assign result_reg_io_enq_valid = io_in_valid; // @[FPU.scala 563:26]
  assign result_reg_io_enq_bits_result = io_in_bits_op == 3'h2 ? {{22'd0}, classifyResult} : _result_T_2; // @[FPU.scala 555:19]
  assign result_reg_io_deq_ready = io_out_ready; // @[FPU.scala 568:26]
endmodule
module RoundingUnit_1(
  input  [2:0]  io_in_rm,
  input  [31:0] io_in_frac,
  input         io_in_sign,
  input         io_in_guard,
  input         io_in_round,
  input         io_in_sticky,
  output [31:0] io_out_fracRounded
);
  wire  inexact = io_in_guard | io_in_round | io_in_sticky; // @[FPU.scala 36:43]
  wire  lsb = io_in_frac[0]; // @[FPU.scala 37:23]
  wire  _roundUp_T_2 = io_in_guard & (io_in_round | io_in_sticky | lsb); // @[FPU.scala 39:25]
  wire  _roundUp_T_4 = inexact & ~io_in_sign; // @[FPU.scala 41:21]
  wire  _roundUp_T_5 = inexact & io_in_sign; // @[FPU.scala 42:21]
  wire  _roundUp_T_9 = 3'h1 == io_in_rm ? 1'h0 : 3'h0 == io_in_rm & _roundUp_T_2; // @[Mux.scala 81:58]
  wire  _roundUp_T_11 = 3'h3 == io_in_rm ? _roundUp_T_4 : _roundUp_T_9; // @[Mux.scala 81:58]
  wire  _roundUp_T_13 = 3'h2 == io_in_rm ? _roundUp_T_5 : _roundUp_T_11; // @[Mux.scala 81:58]
  wire  roundUp = 3'h4 == io_in_rm ? io_in_guard : _roundUp_T_13; // @[Mux.scala 81:58]
  wire [32:0] fracRoundUp = io_in_frac + 32'h1; // @[FPU.scala 45:32]
  assign io_out_fracRounded = roundUp ? fracRoundUp[31:0] : io_in_frac; // @[FPU.scala 47:24]
endmodule
module FPU_F2I(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_op,
  input  [31:0] io_in_bits_a,
  input  [2:0]  io_in_bits_rm,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result
);
  wire [31:0] cls_io_in; // @[FPU.scala 417:19]
  wire  cls_io_isNegInf; // @[FPU.scala 417:19]
  wire  cls_io_isNegNormal; // @[FPU.scala 417:19]
  wire  cls_io_isNegSubnormal; // @[FPU.scala 417:19]
  wire  cls_io_isNegZero; // @[FPU.scala 417:19]
  wire  cls_io_isPosZero; // @[FPU.scala 417:19]
  wire  cls_io_isPosSubnormal; // @[FPU.scala 417:19]
  wire  cls_io_isPosNormal; // @[FPU.scala 417:19]
  wire  cls_io_isPosInf; // @[FPU.scala 417:19]
  wire  cls_io_isSNaN; // @[FPU.scala 417:19]
  wire  cls_io_isQNaN; // @[FPU.scala 417:19]
  wire  cls_io_isNaN; // @[FPU.scala 417:19]
  wire  cls_io_isInf; // @[FPU.scala 417:19]
  wire  cls_io_isInfOrNaN; // @[FPU.scala 417:19]
  wire  cls_io_isSubnormal; // @[FPU.scala 417:19]
  wire  cls_io_isZero; // @[FPU.scala 417:19]
  wire  cls_io_isSubnormalOrZero; // @[FPU.scala 417:19]
  wire [2:0] rounding_io_in_rm; // @[FPU.scala 439:24]
  wire [31:0] rounding_io_in_frac; // @[FPU.scala 439:24]
  wire  rounding_io_in_sign; // @[FPU.scala 439:24]
  wire  rounding_io_in_guard; // @[FPU.scala 439:24]
  wire  rounding_io_in_round; // @[FPU.scala 439:24]
  wire  rounding_io_in_sticky; // @[FPU.scala 439:24]
  wire [31:0] rounding_io_out_fracRounded; // @[FPU.scala 439:24]
  wire  result_reg_clock; // @[FPU.scala 460:24]
  wire  result_reg_reset; // @[FPU.scala 460:24]
  wire  result_reg_io_enq_ready; // @[FPU.scala 460:24]
  wire  result_reg_io_enq_valid; // @[FPU.scala 460:24]
  wire [31:0] result_reg_io_enq_bits_result; // @[FPU.scala 460:24]
  wire  result_reg_io_deq_ready; // @[FPU.scala 460:24]
  wire  result_reg_io_deq_valid; // @[FPU.scala 460:24]
  wire [31:0] result_reg_io_deq_bits_result; // @[FPU.scala 460:24]
  wire [22:0] f32_frac = io_in_bits_a[22:0]; // @[util.scala 46:46]
  wire [7:0] f32_exp = io_in_bits_a[30:23]; // @[util.scala 46:46]
  wire  f32_sign = io_in_bits_a[31]; // @[util.scala 46:46]
  wire [8:0] _exp_T_1 = {1'h0,f32_exp}; // @[util.scala 76:47]
  wire  _frac_T = f32_exp != 8'h0; // @[util.scala 45:33]
  wire [23:0] frac = {_frac_T,f32_frac}; // @[Cat.scala 31:58]
  wire [9:0] exp = {{1{_exp_T_1[8]}},_exp_T_1}; // @[FPU.scala 422:17 423:7]
  wire [9:0] leftShiftAmt = $signed(exp) - 10'sh96; // @[FPU.scala 426:26]
  wire [9:0] _rightShiftAmt_T = $signed(exp) - 10'sh96; // @[FPU.scala 427:43]
  wire [9:0] rightShiftAmt = 10'h0 - _rightShiftAmt_T; // @[FPU.scala 427:23]
  wire  needRightShift = leftShiftAmt[9]; // @[FPU.scala 428:41]
  wire  expOv = $signed(leftShiftAmt) > 10'sh8; // @[FPU.scala 431:28]
  wire [26:0] uintUnrounded_x_ext = {_frac_T,f32_frac,3'h0}; // @[Cat.scala 31:58]
  wire [4:0] uintUnrounded_realShiftAmt = rightShiftAmt > 10'h1a ? 5'h1b : rightShiftAmt[4:0]; // @[util.scala 125:27]
  wire [4:0] _uintUnrounded_mask_T_2 = 5'h1b - uintUnrounded_realShiftAmt; // @[util.scala 129:48]
  wire [26:0] uintUnrounded_mask = 27'h7ffffff >> _uintUnrounded_mask_T_2; // @[util.scala 129:41]
  wire [26:0] uintUnrounded_x_shifted = uintUnrounded_x_ext >> uintUnrounded_realShiftAmt; // @[util.scala 131:24]
  wire [26:0] _uintUnrounded_T_2 = uintUnrounded_mask & uintUnrounded_x_ext; // @[util.scala 132:32]
  wire [26:0] _GEN_0 = {{26'd0}, |_uintUnrounded_T_2}; // @[util.scala 132:23]
  wire [26:0] _uintUnrounded_T_4 = uintUnrounded_x_shifted | _GEN_0; // @[util.scala 132:23]
  wire [38:0] _GEN_1 = {{15'd0}, frac}; // @[FPU.scala 436:15]
  wire [38:0] _uintUnrounded_T_6 = _GEN_1 << leftShiftAmt[3:0]; // @[FPU.scala 436:15]
  wire [34:0] _uintUnrounded_T_8 = {_uintUnrounded_T_6[31:0],3'h0}; // @[Cat.scala 31:58]
  wire [34:0] uintUnrounded = needRightShift ? {{8'd0}, _uintUnrounded_T_4} : _uintUnrounded_T_8; // @[FPU.scala 434:23]
  wire [31:0] _commonResult_T_1 = 32'h0 - rounding_io_out_fracRounded; // @[FPU.scala 448:32]
  wire [31:0] commonResult = f32_sign ? _commonResult_T_1 : rounding_io_out_fracRounded; // @[FPU.scala 448:25]
  wire  _diffSign_T_3 = commonResult[31] ^ f32_sign; // @[FPU.scala 452:22]
  wire  _diffSign_T_4 = io_in_bits_op[0] ? f32_sign : _diffSign_T_3; // @[FPU.scala 450:37]
  wire  diffSign = |rounding_io_out_fracRounded & _diffSign_T_4; // @[FPU.scala 450:31]
  wire [31:0] max32 = {io_in_bits_op[0],31'h7fffffff}; // @[Cat.scala 31:58]
  wire  _min32_T_1 = ~io_in_bits_op[0]; // @[FPU.scala 455:19]
  wire [31:0] min32 = {_min32_T_1,31'h0}; // @[Cat.scala 31:58]
  wire [31:0] specialResult = cls_io_isNaN | ~f32_sign ? max32 : min32; // @[FPU.scala 457:26]
  wire  invalid = cls_io_isNaN | expOv | diffSign; // @[FPU.scala 458:32]
  Classify cls ( // @[FPU.scala 417:19]
    .io_in(cls_io_in),
    .io_isNegInf(cls_io_isNegInf),
    .io_isNegNormal(cls_io_isNegNormal),
    .io_isNegSubnormal(cls_io_isNegSubnormal),
    .io_isNegZero(cls_io_isNegZero),
    .io_isPosZero(cls_io_isPosZero),
    .io_isPosSubnormal(cls_io_isPosSubnormal),
    .io_isPosNormal(cls_io_isPosNormal),
    .io_isPosInf(cls_io_isPosInf),
    .io_isSNaN(cls_io_isSNaN),
    .io_isQNaN(cls_io_isQNaN),
    .io_isNaN(cls_io_isNaN),
    .io_isInf(cls_io_isInf),
    .io_isInfOrNaN(cls_io_isInfOrNaN),
    .io_isSubnormal(cls_io_isSubnormal),
    .io_isZero(cls_io_isZero),
    .io_isSubnormalOrZero(cls_io_isSubnormalOrZero)
  );
  RoundingUnit_1 rounding ( // @[FPU.scala 439:24]
    .io_in_rm(rounding_io_in_rm),
    .io_in_frac(rounding_io_in_frac),
    .io_in_sign(rounding_io_in_sign),
    .io_in_guard(rounding_io_in_guard),
    .io_in_round(rounding_io_in_round),
    .io_in_sticky(rounding_io_in_sticky),
    .io_out_fracRounded(rounding_io_out_fracRounded)
  );
  Queue_5 result_reg ( // @[FPU.scala 460:24]
    .clock(result_reg_clock),
    .reset(result_reg_reset),
    .io_enq_ready(result_reg_io_enq_ready),
    .io_enq_valid(result_reg_io_enq_valid),
    .io_enq_bits_result(result_reg_io_enq_bits_result),
    .io_deq_ready(result_reg_io_deq_ready),
    .io_deq_valid(result_reg_io_deq_valid),
    .io_deq_bits_result(result_reg_io_deq_bits_result)
  );
  assign io_in_ready = result_reg_io_enq_ready; // @[FPU.scala 468:14]
  assign io_out_valid = result_reg_io_deq_valid; // @[FPU.scala 470:16]
  assign io_out_bits_result = result_reg_io_deq_bits_result; // @[FPU.scala 471:14]
  assign cls_io_in = io_in_bits_a; // @[FPU.scala 418:13]
  assign rounding_io_in_rm = io_in_bits_rm; // @[FPU.scala 440:21]
  assign rounding_io_in_frac = uintUnrounded[34:3]; // @[FPU.scala 442:44]
  assign rounding_io_in_sign = io_in_bits_a[31]; // @[util.scala 46:46]
  assign rounding_io_in_guard = uintUnrounded[2]; // @[FPU.scala 443:54]
  assign rounding_io_in_round = uintUnrounded[1]; // @[FPU.scala 444:54]
  assign rounding_io_in_sticky = uintUnrounded[0]; // @[FPU.scala 445:46]
  assign result_reg_clock = clock;
  assign result_reg_reset = reset;
  assign result_reg_io_enq_valid = io_in_valid; // @[FPU.scala 467:26]
  assign result_reg_io_enq_bits_result = invalid ? specialResult : commonResult; // @[FPU.scala 461:39]
  assign result_reg_io_deq_ready = io_out_ready; // @[FPU.scala 472:26]
endmodule
module RoundingUnit_2(
  input  [2:0]  io_in_rm,
  input  [22:0] io_in_frac,
  input         io_in_sign,
  input         io_in_guard,
  input         io_in_round,
  input         io_in_sticky,
  output [22:0] io_out_fracRounded,
  output        io_out_fracCout
);
  wire  inexact = io_in_guard | io_in_round | io_in_sticky; // @[FPU.scala 36:43]
  wire  lsb = io_in_frac[0]; // @[FPU.scala 37:23]
  wire  _roundUp_T_2 = io_in_guard & (io_in_round | io_in_sticky | lsb); // @[FPU.scala 39:25]
  wire  _roundUp_T_4 = inexact & ~io_in_sign; // @[FPU.scala 41:21]
  wire  _roundUp_T_5 = inexact & io_in_sign; // @[FPU.scala 42:21]
  wire  _roundUp_T_9 = 3'h1 == io_in_rm ? 1'h0 : 3'h0 == io_in_rm & _roundUp_T_2; // @[Mux.scala 81:58]
  wire  _roundUp_T_11 = 3'h3 == io_in_rm ? _roundUp_T_4 : _roundUp_T_9; // @[Mux.scala 81:58]
  wire  _roundUp_T_13 = 3'h2 == io_in_rm ? _roundUp_T_5 : _roundUp_T_11; // @[Mux.scala 81:58]
  wire  roundUp = 3'h4 == io_in_rm ? io_in_guard : _roundUp_T_13; // @[Mux.scala 81:58]
  wire [23:0] fracRoundUp = io_in_frac + 23'h1; // @[FPU.scala 45:32]
  wire  cout = fracRoundUp[23]; // @[FPU.scala 46:25]
  assign io_out_fracRounded = roundUp ? fracRoundUp[22:0] : io_in_frac; // @[FPU.scala 47:24]
  assign io_out_fracCout = cout & roundUp; // @[FPU.scala 50:27]
endmodule
module FPU_I2F(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_op,
  input  [31:0] io_in_bits_a,
  input  [2:0]  io_in_bits_rm,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result
);
  wire [2:0] roundingUnit_io_in_rm; // @[FPU.scala 500:28]
  wire [22:0] roundingUnit_io_in_frac; // @[FPU.scala 500:28]
  wire  roundingUnit_io_in_sign; // @[FPU.scala 500:28]
  wire  roundingUnit_io_in_guard; // @[FPU.scala 500:28]
  wire  roundingUnit_io_in_round; // @[FPU.scala 500:28]
  wire  roundingUnit_io_in_sticky; // @[FPU.scala 500:28]
  wire [22:0] roundingUnit_io_out_fracRounded; // @[FPU.scala 500:28]
  wire  roundingUnit_io_out_fracCout; // @[FPU.scala 500:28]
  wire  result_reg_clock; // @[FPU.scala 517:24]
  wire  result_reg_reset; // @[FPU.scala 517:24]
  wire  result_reg_io_enq_ready; // @[FPU.scala 517:24]
  wire  result_reg_io_enq_valid; // @[FPU.scala 517:24]
  wire [31:0] result_reg_io_enq_bits_result; // @[FPU.scala 517:24]
  wire  result_reg_io_deq_ready; // @[FPU.scala 517:24]
  wire  result_reg_io_deq_valid; // @[FPU.scala 517:24]
  wire [31:0] result_reg_io_deq_bits_result; // @[FPU.scala 517:24]
  wire [31:0] aNeg = ~io_in_bits_a; // @[FPU.scala 479:15]
  wire [31:0] aComp = aNeg + 32'h1; // @[FPU.scala 480:20]
  wire  aSign = io_in_bits_op[0] ? 1'h0 : io_in_bits_a[31]; // @[FPU.scala 481:18]
  wire [4:0] _leadingZerosComp_T_32 = aComp[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_33 = aComp[2] ? 5'h1d : _leadingZerosComp_T_32; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_34 = aComp[3] ? 5'h1c : _leadingZerosComp_T_33; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_35 = aComp[4] ? 5'h1b : _leadingZerosComp_T_34; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_36 = aComp[5] ? 5'h1a : _leadingZerosComp_T_35; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_37 = aComp[6] ? 5'h19 : _leadingZerosComp_T_36; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_38 = aComp[7] ? 5'h18 : _leadingZerosComp_T_37; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_39 = aComp[8] ? 5'h17 : _leadingZerosComp_T_38; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_40 = aComp[9] ? 5'h16 : _leadingZerosComp_T_39; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_41 = aComp[10] ? 5'h15 : _leadingZerosComp_T_40; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_42 = aComp[11] ? 5'h14 : _leadingZerosComp_T_41; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_43 = aComp[12] ? 5'h13 : _leadingZerosComp_T_42; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_44 = aComp[13] ? 5'h12 : _leadingZerosComp_T_43; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_45 = aComp[14] ? 5'h11 : _leadingZerosComp_T_44; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_46 = aComp[15] ? 5'h10 : _leadingZerosComp_T_45; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_47 = aComp[16] ? 5'hf : _leadingZerosComp_T_46; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_48 = aComp[17] ? 5'he : _leadingZerosComp_T_47; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_49 = aComp[18] ? 5'hd : _leadingZerosComp_T_48; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_50 = aComp[19] ? 5'hc : _leadingZerosComp_T_49; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_51 = aComp[20] ? 5'hb : _leadingZerosComp_T_50; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_52 = aComp[21] ? 5'ha : _leadingZerosComp_T_51; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_53 = aComp[22] ? 5'h9 : _leadingZerosComp_T_52; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_54 = aComp[23] ? 5'h8 : _leadingZerosComp_T_53; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_55 = aComp[24] ? 5'h7 : _leadingZerosComp_T_54; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_56 = aComp[25] ? 5'h6 : _leadingZerosComp_T_55; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_57 = aComp[26] ? 5'h5 : _leadingZerosComp_T_56; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_58 = aComp[27] ? 5'h4 : _leadingZerosComp_T_57; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_59 = aComp[28] ? 5'h3 : _leadingZerosComp_T_58; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_60 = aComp[29] ? 5'h2 : _leadingZerosComp_T_59; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosComp_T_61 = aComp[30] ? 5'h1 : _leadingZerosComp_T_60; // @[Mux.scala 47:70]
  wire [4:0] leadingZerosComp = aComp[31] ? 5'h0 : _leadingZerosComp_T_61; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_32 = aNeg[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_33 = aNeg[2] ? 5'h1d : _leadingZerosNeg_T_32; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_34 = aNeg[3] ? 5'h1c : _leadingZerosNeg_T_33; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_35 = aNeg[4] ? 5'h1b : _leadingZerosNeg_T_34; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_36 = aNeg[5] ? 5'h1a : _leadingZerosNeg_T_35; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_37 = aNeg[6] ? 5'h19 : _leadingZerosNeg_T_36; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_38 = aNeg[7] ? 5'h18 : _leadingZerosNeg_T_37; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_39 = aNeg[8] ? 5'h17 : _leadingZerosNeg_T_38; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_40 = aNeg[9] ? 5'h16 : _leadingZerosNeg_T_39; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_41 = aNeg[10] ? 5'h15 : _leadingZerosNeg_T_40; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_42 = aNeg[11] ? 5'h14 : _leadingZerosNeg_T_41; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_43 = aNeg[12] ? 5'h13 : _leadingZerosNeg_T_42; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_44 = aNeg[13] ? 5'h12 : _leadingZerosNeg_T_43; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_45 = aNeg[14] ? 5'h11 : _leadingZerosNeg_T_44; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_46 = aNeg[15] ? 5'h10 : _leadingZerosNeg_T_45; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_47 = aNeg[16] ? 5'hf : _leadingZerosNeg_T_46; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_48 = aNeg[17] ? 5'he : _leadingZerosNeg_T_47; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_49 = aNeg[18] ? 5'hd : _leadingZerosNeg_T_48; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_50 = aNeg[19] ? 5'hc : _leadingZerosNeg_T_49; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_51 = aNeg[20] ? 5'hb : _leadingZerosNeg_T_50; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_52 = aNeg[21] ? 5'ha : _leadingZerosNeg_T_51; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_53 = aNeg[22] ? 5'h9 : _leadingZerosNeg_T_52; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_54 = aNeg[23] ? 5'h8 : _leadingZerosNeg_T_53; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_55 = aNeg[24] ? 5'h7 : _leadingZerosNeg_T_54; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_56 = aNeg[25] ? 5'h6 : _leadingZerosNeg_T_55; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_57 = aNeg[26] ? 5'h5 : _leadingZerosNeg_T_56; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_58 = aNeg[27] ? 5'h4 : _leadingZerosNeg_T_57; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_59 = aNeg[28] ? 5'h3 : _leadingZerosNeg_T_58; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_60 = aNeg[29] ? 5'h2 : _leadingZerosNeg_T_59; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosNeg_T_61 = aNeg[30] ? 5'h1 : _leadingZerosNeg_T_60; // @[Mux.scala 47:70]
  wire [4:0] leadingZerosNeg = aNeg[31] ? 5'h0 : _leadingZerosNeg_T_61; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_32 = io_in_bits_a[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_33 = io_in_bits_a[2] ? 5'h1d : _leadingZerosPos_T_32; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_34 = io_in_bits_a[3] ? 5'h1c : _leadingZerosPos_T_33; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_35 = io_in_bits_a[4] ? 5'h1b : _leadingZerosPos_T_34; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_36 = io_in_bits_a[5] ? 5'h1a : _leadingZerosPos_T_35; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_37 = io_in_bits_a[6] ? 5'h19 : _leadingZerosPos_T_36; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_38 = io_in_bits_a[7] ? 5'h18 : _leadingZerosPos_T_37; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_39 = io_in_bits_a[8] ? 5'h17 : _leadingZerosPos_T_38; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_40 = io_in_bits_a[9] ? 5'h16 : _leadingZerosPos_T_39; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_41 = io_in_bits_a[10] ? 5'h15 : _leadingZerosPos_T_40; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_42 = io_in_bits_a[11] ? 5'h14 : _leadingZerosPos_T_41; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_43 = io_in_bits_a[12] ? 5'h13 : _leadingZerosPos_T_42; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_44 = io_in_bits_a[13] ? 5'h12 : _leadingZerosPos_T_43; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_45 = io_in_bits_a[14] ? 5'h11 : _leadingZerosPos_T_44; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_46 = io_in_bits_a[15] ? 5'h10 : _leadingZerosPos_T_45; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_47 = io_in_bits_a[16] ? 5'hf : _leadingZerosPos_T_46; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_48 = io_in_bits_a[17] ? 5'he : _leadingZerosPos_T_47; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_49 = io_in_bits_a[18] ? 5'hd : _leadingZerosPos_T_48; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_50 = io_in_bits_a[19] ? 5'hc : _leadingZerosPos_T_49; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_51 = io_in_bits_a[20] ? 5'hb : _leadingZerosPos_T_50; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_52 = io_in_bits_a[21] ? 5'ha : _leadingZerosPos_T_51; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_53 = io_in_bits_a[22] ? 5'h9 : _leadingZerosPos_T_52; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_54 = io_in_bits_a[23] ? 5'h8 : _leadingZerosPos_T_53; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_55 = io_in_bits_a[24] ? 5'h7 : _leadingZerosPos_T_54; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_56 = io_in_bits_a[25] ? 5'h6 : _leadingZerosPos_T_55; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_57 = io_in_bits_a[26] ? 5'h5 : _leadingZerosPos_T_56; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_58 = io_in_bits_a[27] ? 5'h4 : _leadingZerosPos_T_57; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_59 = io_in_bits_a[28] ? 5'h3 : _leadingZerosPos_T_58; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_60 = io_in_bits_a[29] ? 5'h2 : _leadingZerosPos_T_59; // @[Mux.scala 47:70]
  wire [4:0] _leadingZerosPos_T_61 = io_in_bits_a[30] ? 5'h1 : _leadingZerosPos_T_60; // @[Mux.scala 47:70]
  wire [4:0] leadingZerosPos = io_in_bits_a[31] ? 5'h0 : _leadingZerosPos_T_61; // @[Mux.scala 47:70]
  wire [31:0] aVal = aSign ? aComp : io_in_bits_a; // @[FPU.scala 487:17]
  wire [4:0] leadingZeros = aSign ? leadingZerosNeg : leadingZerosPos; // @[FPU.scala 488:25]
  wire [7:0] _GEN_0 = {{3'd0}, leadingZeros}; // @[FPU.scala 490:54]
  wire [7:0] expUnrounded = 8'h9e - _GEN_0; // @[FPU.scala 490:54]
  wire  leadingZeroHasError = aSign & leadingZerosComp != leadingZerosNeg; // @[FPU.scala 491:35]
  wire [62:0] _GEN_3 = {{31'd0}, aVal}; // @[FPU.scala 492:23]
  wire [62:0] _aShifted_T = _GEN_3 << leadingZeros; // @[FPU.scala 492:23]
  wire [31:0] aShifted = _aShifted_T[31:0]; // @[FPU.scala 492:38]
  wire [30:0] aShiftedFix = leadingZeroHasError ? aShifted[31:1] : aShifted[30:0]; // @[FPU.scala 494:24]
  wire [7:0] _GEN_1 = {{7'd0}, roundingUnit_io_out_fracCout}; // @[FPU.scala 509:33]
  wire [7:0] _expRounded_T_1 = expUnrounded + _GEN_1; // @[FPU.scala 509:33]
  wire [7:0] _GEN_2 = {{7'd0}, leadingZeroHasError}; // @[FPU.scala 509:64]
  wire [7:0] expRounded = _expRounded_T_1 + _GEN_2; // @[FPU.scala 509:64]
  wire [22:0] _resF_T_1 = roundingUnit_io_out_fracRounded; // @[FPU.scala 514:16]
  wire [31:0] resF = {aSign,expRounded,_resF_T_1}; // @[Cat.scala 31:58]
  RoundingUnit_2 roundingUnit ( // @[FPU.scala 500:28]
    .io_in_rm(roundingUnit_io_in_rm),
    .io_in_frac(roundingUnit_io_in_frac),
    .io_in_sign(roundingUnit_io_in_sign),
    .io_in_guard(roundingUnit_io_in_guard),
    .io_in_round(roundingUnit_io_in_round),
    .io_in_sticky(roundingUnit_io_in_sticky),
    .io_out_fracRounded(roundingUnit_io_out_fracRounded),
    .io_out_fracCout(roundingUnit_io_out_fracCout)
  );
  Queue_5 result_reg ( // @[FPU.scala 517:24]
    .clock(result_reg_clock),
    .reset(result_reg_reset),
    .io_enq_ready(result_reg_io_enq_ready),
    .io_enq_valid(result_reg_io_enq_valid),
    .io_enq_bits_result(result_reg_io_enq_bits_result),
    .io_deq_ready(result_reg_io_deq_ready),
    .io_deq_valid(result_reg_io_deq_valid),
    .io_deq_bits_result(result_reg_io_deq_bits_result)
  );
  assign io_in_ready = result_reg_io_enq_ready; // @[FPU.scala 525:14]
  assign io_out_valid = result_reg_io_deq_valid; // @[FPU.scala 527:16]
  assign io_out_bits_result = result_reg_io_deq_bits_result; // @[FPU.scala 528:14]
  assign roundingUnit_io_in_rm = io_in_bits_rm; // @[FPU.scala 501:25]
  assign roundingUnit_io_in_frac = aShiftedFix[30:8]; // @[FPU.scala 495:26]
  assign roundingUnit_io_in_sign = io_in_bits_op[0] ? 1'h0 : io_in_bits_a[31]; // @[FPU.scala 481:18]
  assign roundingUnit_io_in_guard = aShiftedFix[7]; // @[FPU.scala 496:22]
  assign roundingUnit_io_in_round = aShiftedFix[6]; // @[FPU.scala 497:22]
  assign roundingUnit_io_in_sticky = |aShiftedFix[5:0]; // @[FPU.scala 498:35]
  assign result_reg_clock = clock;
  assign result_reg_reset = reset;
  assign result_reg_io_enq_valid = io_in_valid; // @[FPU.scala 524:26]
  assign result_reg_io_enq_bits_result = io_in_bits_a == 32'h0 ? 32'h0 : resF; // @[FPU.scala 518:39]
  assign result_reg_io_deq_ready = io_out_ready; // @[FPU.scala 529:26]
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_result,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_result,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_result,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_result,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [31:0] io_in_4_bits_result,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result,
  output [2:0]  io_chosen
);
  wire [2:0] _GEN_0 = io_in_3_valid ? 3'h3 : 3'h4; // @[Arbiter.scala 138:13 141:26 142:17]
  wire [31:0] _GEN_6 = io_in_3_valid ? io_in_3_bits_result : io_in_4_bits_result; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [2:0] _GEN_7 = io_in_2_valid ? 3'h2 : _GEN_0; // @[Arbiter.scala 141:26 142:17]
  wire [31:0] _GEN_13 = io_in_2_valid ? io_in_2_bits_result : _GEN_6; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_14 = io_in_1_valid ? 3'h1 : _GEN_7; // @[Arbiter.scala 141:26 142:17]
  wire [31:0] _GEN_20 = io_in_1_valid ? io_in_1_bits_result : _GEN_13; // @[Arbiter.scala 141:26 143:19]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 46:78]
  wire  grant_3 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 46:78]
  wire  grant_4 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid); // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_2_ready = grant_2 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_3_ready = grant_3 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_4_ready = grant_4 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_4 | io_in_4_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_result = io_in_0_valid ? io_in_0_bits_result : _GEN_20; // @[Arbiter.scala 141:26 143:19]
  assign io_chosen = io_in_0_valid ? 3'h0 : _GEN_14; // @[Arbiter.scala 141:26 142:17]
endmodule
module ScalarFPU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [5:0]  io_in_bits_fpuop,
  input  [31:0] io_in_bits_a,
  input  [31:0] io_in_bits_b,
  input  [31:0] io_in_bits_c,
  input  [2:0]  io_in_bits_rm,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result,
  output [2:0]  io_select
);
  wire  FPU_FMA_clock; // @[FPU.scala 587:11]
  wire  FPU_FMA_reset; // @[FPU.scala 587:11]
  wire  FPU_FMA_io_in_ready; // @[FPU.scala 587:11]
  wire  FPU_FMA_io_in_valid; // @[FPU.scala 587:11]
  wire [2:0] FPU_FMA_io_in_bits_op; // @[FPU.scala 587:11]
  wire [31:0] FPU_FMA_io_in_bits_a; // @[FPU.scala 587:11]
  wire [31:0] FPU_FMA_io_in_bits_b; // @[FPU.scala 587:11]
  wire [31:0] FPU_FMA_io_in_bits_c; // @[FPU.scala 587:11]
  wire [2:0] FPU_FMA_io_in_bits_rm; // @[FPU.scala 587:11]
  wire  FPU_FMA_io_out_ready; // @[FPU.scala 587:11]
  wire  FPU_FMA_io_out_valid; // @[FPU.scala 587:11]
  wire [31:0] FPU_FMA_io_out_bits_result; // @[FPU.scala 587:11]
  wire  FPU_CMP_clock; // @[FPU.scala 588:11]
  wire  FPU_CMP_reset; // @[FPU.scala 588:11]
  wire  FPU_CMP_io_in_ready; // @[FPU.scala 588:11]
  wire  FPU_CMP_io_in_valid; // @[FPU.scala 588:11]
  wire [2:0] FPU_CMP_io_in_bits_op; // @[FPU.scala 588:11]
  wire [31:0] FPU_CMP_io_in_bits_a; // @[FPU.scala 588:11]
  wire [31:0] FPU_CMP_io_in_bits_b; // @[FPU.scala 588:11]
  wire  FPU_CMP_io_out_ready; // @[FPU.scala 588:11]
  wire  FPU_CMP_io_out_valid; // @[FPU.scala 588:11]
  wire [31:0] FPU_CMP_io_out_bits_result; // @[FPU.scala 588:11]
  wire  FPU_FMV_clock; // @[FPU.scala 589:11]
  wire  FPU_FMV_reset; // @[FPU.scala 589:11]
  wire  FPU_FMV_io_in_ready; // @[FPU.scala 589:11]
  wire  FPU_FMV_io_in_valid; // @[FPU.scala 589:11]
  wire [2:0] FPU_FMV_io_in_bits_op; // @[FPU.scala 589:11]
  wire [31:0] FPU_FMV_io_in_bits_a; // @[FPU.scala 589:11]
  wire [31:0] FPU_FMV_io_in_bits_b; // @[FPU.scala 589:11]
  wire  FPU_FMV_io_out_ready; // @[FPU.scala 589:11]
  wire  FPU_FMV_io_out_valid; // @[FPU.scala 589:11]
  wire [31:0] FPU_FMV_io_out_bits_result; // @[FPU.scala 589:11]
  wire  FPU_F2I_clock; // @[FPU.scala 590:11]
  wire  FPU_F2I_reset; // @[FPU.scala 590:11]
  wire  FPU_F2I_io_in_ready; // @[FPU.scala 590:11]
  wire  FPU_F2I_io_in_valid; // @[FPU.scala 590:11]
  wire [2:0] FPU_F2I_io_in_bits_op; // @[FPU.scala 590:11]
  wire [31:0] FPU_F2I_io_in_bits_a; // @[FPU.scala 590:11]
  wire [2:0] FPU_F2I_io_in_bits_rm; // @[FPU.scala 590:11]
  wire  FPU_F2I_io_out_ready; // @[FPU.scala 590:11]
  wire  FPU_F2I_io_out_valid; // @[FPU.scala 590:11]
  wire [31:0] FPU_F2I_io_out_bits_result; // @[FPU.scala 590:11]
  wire  FPU_I2F_clock; // @[FPU.scala 591:11]
  wire  FPU_I2F_reset; // @[FPU.scala 591:11]
  wire  FPU_I2F_io_in_ready; // @[FPU.scala 591:11]
  wire  FPU_I2F_io_in_valid; // @[FPU.scala 591:11]
  wire [2:0] FPU_I2F_io_in_bits_op; // @[FPU.scala 591:11]
  wire [31:0] FPU_I2F_io_in_bits_a; // @[FPU.scala 591:11]
  wire [2:0] FPU_I2F_io_in_bits_rm; // @[FPU.scala 591:11]
  wire  FPU_I2F_io_out_ready; // @[FPU.scala 591:11]
  wire  FPU_I2F_io_out_valid; // @[FPU.scala 591:11]
  wire [31:0] FPU_I2F_io_out_bits_result; // @[FPU.scala 591:11]
  wire  outArbiter_io_in_0_ready; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_0_valid; // @[FPU.scala 613:26]
  wire [31:0] outArbiter_io_in_0_bits_result; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_1_ready; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_1_valid; // @[FPU.scala 613:26]
  wire [31:0] outArbiter_io_in_1_bits_result; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_2_ready; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_2_valid; // @[FPU.scala 613:26]
  wire [31:0] outArbiter_io_in_2_bits_result; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_3_ready; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_3_valid; // @[FPU.scala 613:26]
  wire [31:0] outArbiter_io_in_3_bits_result; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_4_ready; // @[FPU.scala 613:26]
  wire  outArbiter_io_in_4_valid; // @[FPU.scala 613:26]
  wire [31:0] outArbiter_io_in_4_bits_result; // @[FPU.scala 613:26]
  wire  outArbiter_io_out_ready; // @[FPU.scala 613:26]
  wire  outArbiter_io_out_valid; // @[FPU.scala 613:26]
  wire [31:0] outArbiter_io_out_bits_result; // @[FPU.scala 613:26]
  wire [2:0] outArbiter_io_chosen; // @[FPU.scala 613:26]
  wire [2:0] fu = io_in_bits_fpuop[5:3]; // @[FPU.scala 584:28]
  wire [2:0] op = io_in_bits_fpuop[2:0]; // @[FPU.scala 585:28]
  wire  _T = 3'h0 == fu; // @[FPU.scala 595:41]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & FPU_FMA_io_in_ready; // @[FPU.scala 593:14 601:{21,33}]
  wire  _T_14 = 3'h1 == fu; // @[FPU.scala 595:41]
  wire  _GEN_1 = _T_14 ? FPU_CMP_io_in_ready : _GEN_0; // @[FPU.scala 601:{21,33}]
  wire  _T_28 = 3'h2 == fu; // @[FPU.scala 595:41]
  wire  _GEN_2 = _T_28 ? FPU_FMV_io_in_ready : _GEN_1; // @[FPU.scala 601:{21,33}]
  wire  _T_42 = 3'h3 == fu; // @[FPU.scala 595:41]
  wire  _GEN_3 = _T_42 ? FPU_F2I_io_in_ready : _GEN_2; // @[FPU.scala 601:{21,33}]
  wire  _T_56 = 3'h4 == fu; // @[FPU.scala 595:41]
  FPU_FMA FPU_FMA ( // @[FPU.scala 587:11]
    .clock(FPU_FMA_clock),
    .reset(FPU_FMA_reset),
    .io_in_ready(FPU_FMA_io_in_ready),
    .io_in_valid(FPU_FMA_io_in_valid),
    .io_in_bits_op(FPU_FMA_io_in_bits_op),
    .io_in_bits_a(FPU_FMA_io_in_bits_a),
    .io_in_bits_b(FPU_FMA_io_in_bits_b),
    .io_in_bits_c(FPU_FMA_io_in_bits_c),
    .io_in_bits_rm(FPU_FMA_io_in_bits_rm),
    .io_out_ready(FPU_FMA_io_out_ready),
    .io_out_valid(FPU_FMA_io_out_valid),
    .io_out_bits_result(FPU_FMA_io_out_bits_result)
  );
  FPU_CMP FPU_CMP ( // @[FPU.scala 588:11]
    .clock(FPU_CMP_clock),
    .reset(FPU_CMP_reset),
    .io_in_ready(FPU_CMP_io_in_ready),
    .io_in_valid(FPU_CMP_io_in_valid),
    .io_in_bits_op(FPU_CMP_io_in_bits_op),
    .io_in_bits_a(FPU_CMP_io_in_bits_a),
    .io_in_bits_b(FPU_CMP_io_in_bits_b),
    .io_out_ready(FPU_CMP_io_out_ready),
    .io_out_valid(FPU_CMP_io_out_valid),
    .io_out_bits_result(FPU_CMP_io_out_bits_result)
  );
  FPU_FMV FPU_FMV ( // @[FPU.scala 589:11]
    .clock(FPU_FMV_clock),
    .reset(FPU_FMV_reset),
    .io_in_ready(FPU_FMV_io_in_ready),
    .io_in_valid(FPU_FMV_io_in_valid),
    .io_in_bits_op(FPU_FMV_io_in_bits_op),
    .io_in_bits_a(FPU_FMV_io_in_bits_a),
    .io_in_bits_b(FPU_FMV_io_in_bits_b),
    .io_out_ready(FPU_FMV_io_out_ready),
    .io_out_valid(FPU_FMV_io_out_valid),
    .io_out_bits_result(FPU_FMV_io_out_bits_result)
  );
  FPU_F2I FPU_F2I ( // @[FPU.scala 590:11]
    .clock(FPU_F2I_clock),
    .reset(FPU_F2I_reset),
    .io_in_ready(FPU_F2I_io_in_ready),
    .io_in_valid(FPU_F2I_io_in_valid),
    .io_in_bits_op(FPU_F2I_io_in_bits_op),
    .io_in_bits_a(FPU_F2I_io_in_bits_a),
    .io_in_bits_rm(FPU_F2I_io_in_bits_rm),
    .io_out_ready(FPU_F2I_io_out_ready),
    .io_out_valid(FPU_F2I_io_out_valid),
    .io_out_bits_result(FPU_F2I_io_out_bits_result)
  );
  FPU_I2F FPU_I2F ( // @[FPU.scala 591:11]
    .clock(FPU_I2F_clock),
    .reset(FPU_I2F_reset),
    .io_in_ready(FPU_I2F_io_in_ready),
    .io_in_valid(FPU_I2F_io_in_valid),
    .io_in_bits_op(FPU_I2F_io_in_bits_op),
    .io_in_bits_a(FPU_I2F_io_in_bits_a),
    .io_in_bits_rm(FPU_I2F_io_in_bits_rm),
    .io_out_ready(FPU_I2F_io_out_ready),
    .io_out_valid(FPU_I2F_io_out_valid),
    .io_out_bits_result(FPU_I2F_io_out_bits_result)
  );
  Arbiter outArbiter ( // @[FPU.scala 613:26]
    .io_in_0_ready(outArbiter_io_in_0_ready),
    .io_in_0_valid(outArbiter_io_in_0_valid),
    .io_in_0_bits_result(outArbiter_io_in_0_bits_result),
    .io_in_1_ready(outArbiter_io_in_1_ready),
    .io_in_1_valid(outArbiter_io_in_1_valid),
    .io_in_1_bits_result(outArbiter_io_in_1_bits_result),
    .io_in_2_ready(outArbiter_io_in_2_ready),
    .io_in_2_valid(outArbiter_io_in_2_valid),
    .io_in_2_bits_result(outArbiter_io_in_2_bits_result),
    .io_in_3_ready(outArbiter_io_in_3_ready),
    .io_in_3_valid(outArbiter_io_in_3_valid),
    .io_in_3_bits_result(outArbiter_io_in_3_bits_result),
    .io_in_4_ready(outArbiter_io_in_4_ready),
    .io_in_4_valid(outArbiter_io_in_4_valid),
    .io_in_4_bits_result(outArbiter_io_in_4_bits_result),
    .io_out_ready(outArbiter_io_out_ready),
    .io_out_valid(outArbiter_io_out_valid),
    .io_out_bits_result(outArbiter_io_out_bits_result),
    .io_chosen(outArbiter_io_chosen)
  );
  assign io_in_ready = _T_56 ? FPU_I2F_io_in_ready : _GEN_3; // @[FPU.scala 601:{21,33}]
  assign io_out_valid = outArbiter_io_out_valid; // @[FPU.scala 619:10]
  assign io_out_bits_result = outArbiter_io_out_bits_result; // @[FPU.scala 619:10]
  assign io_select = outArbiter_io_chosen; // @[FPU.scala 620:12]
  assign FPU_FMA_clock = clock;
  assign FPU_FMA_reset = reset;
  assign FPU_FMA_io_in_valid = _T_10 & _T; // @[FPU.scala 600:45]
  assign FPU_FMA_io_in_bits_op = 3'h0 == fu ? op : 3'h0; // @[FPU.scala 595:35]
  assign FPU_FMA_io_in_bits_a = _T ? io_in_bits_a : 32'h0; // @[FPU.scala 597:35]
  assign FPU_FMA_io_in_bits_b = _T ? io_in_bits_b : 32'h0; // @[FPU.scala 598:35]
  assign FPU_FMA_io_in_bits_c = _T ? io_in_bits_c : 32'h0; // @[FPU.scala 599:35]
  assign FPU_FMA_io_in_bits_rm = _T ? io_in_bits_rm : 3'h0; // @[FPU.scala 596:35]
  assign FPU_FMA_io_out_ready = outArbiter_io_in_0_ready; // @[FPU.scala 617:27]
  assign FPU_CMP_clock = clock;
  assign FPU_CMP_reset = reset;
  assign FPU_CMP_io_in_valid = _T_10 & _T_14; // @[FPU.scala 600:45]
  assign FPU_CMP_io_in_bits_op = 3'h1 == fu ? op : 3'h0; // @[FPU.scala 595:35]
  assign FPU_CMP_io_in_bits_a = _T_14 ? io_in_bits_a : 32'h0; // @[FPU.scala 597:35]
  assign FPU_CMP_io_in_bits_b = _T_14 ? io_in_bits_b : 32'h0; // @[FPU.scala 598:35]
  assign FPU_CMP_io_out_ready = outArbiter_io_in_1_ready; // @[FPU.scala 617:27]
  assign FPU_FMV_clock = clock;
  assign FPU_FMV_reset = reset;
  assign FPU_FMV_io_in_valid = _T_10 & _T_28; // @[FPU.scala 600:45]
  assign FPU_FMV_io_in_bits_op = 3'h2 == fu ? op : 3'h0; // @[FPU.scala 595:35]
  assign FPU_FMV_io_in_bits_a = _T_28 ? io_in_bits_a : 32'h0; // @[FPU.scala 597:35]
  assign FPU_FMV_io_in_bits_b = _T_28 ? io_in_bits_b : 32'h0; // @[FPU.scala 598:35]
  assign FPU_FMV_io_out_ready = outArbiter_io_in_2_ready; // @[FPU.scala 617:27]
  assign FPU_F2I_clock = clock;
  assign FPU_F2I_reset = reset;
  assign FPU_F2I_io_in_valid = _T_10 & _T_42; // @[FPU.scala 600:45]
  assign FPU_F2I_io_in_bits_op = 3'h3 == fu ? op : 3'h0; // @[FPU.scala 595:35]
  assign FPU_F2I_io_in_bits_a = _T_42 ? io_in_bits_a : 32'h0; // @[FPU.scala 597:35]
  assign FPU_F2I_io_in_bits_rm = _T_42 ? io_in_bits_rm : 3'h0; // @[FPU.scala 596:35]
  assign FPU_F2I_io_out_ready = outArbiter_io_in_3_ready; // @[FPU.scala 617:27]
  assign FPU_I2F_clock = clock;
  assign FPU_I2F_reset = reset;
  assign FPU_I2F_io_in_valid = _T_10 & _T_56; // @[FPU.scala 600:45]
  assign FPU_I2F_io_in_bits_op = 3'h4 == fu ? op : 3'h0; // @[FPU.scala 595:35]
  assign FPU_I2F_io_in_bits_a = _T_56 ? io_in_bits_a : 32'h0; // @[FPU.scala 597:35]
  assign FPU_I2F_io_in_bits_rm = _T_56 ? io_in_bits_rm : 3'h0; // @[FPU.scala 596:35]
  assign FPU_I2F_io_out_ready = outArbiter_io_in_4_ready; // @[FPU.scala 617:27]
  assign outArbiter_io_in_0_valid = FPU_FMA_io_out_valid; // @[FPU.scala 617:27]
  assign outArbiter_io_in_0_bits_result = FPU_FMA_io_out_bits_result; // @[FPU.scala 617:27]
  assign outArbiter_io_in_1_valid = FPU_CMP_io_out_valid; // @[FPU.scala 617:27]
  assign outArbiter_io_in_1_bits_result = FPU_CMP_io_out_bits_result; // @[FPU.scala 617:27]
  assign outArbiter_io_in_2_valid = FPU_FMV_io_out_valid; // @[FPU.scala 617:27]
  assign outArbiter_io_in_2_bits_result = FPU_FMV_io_out_bits_result; // @[FPU.scala 617:27]
  assign outArbiter_io_in_3_valid = FPU_F2I_io_out_valid; // @[FPU.scala 617:27]
  assign outArbiter_io_in_3_bits_result = FPU_F2I_io_out_bits_result; // @[FPU.scala 617:27]
  assign outArbiter_io_in_4_valid = FPU_I2F_io_out_valid; // @[FPU.scala 617:27]
  assign outArbiter_io_in_4_bits_result = FPU_I2F_io_out_bits_result; // @[FPU.scala 617:27]
  assign outArbiter_io_out_ready = io_out_ready; // @[FPU.scala 619:10]
endmodule
module Queue_39(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits_ctrl_wid,
  input  [4:0] io_enq_bits_ctrl_reg_idxw,
  input        io_enq_bits_ctrl_wfd,
  input        io_enq_bits_ctrl_wxd,
  input        io_enq_bits_mask_0,
  input        io_enq_bits_mask_1,
  input        io_enq_bits_mask_2,
  input        io_enq_bits_mask_3,
  input        io_enq_bits_mask_4,
  input        io_enq_bits_mask_5,
  input        io_enq_bits_mask_6,
  input        io_enq_bits_mask_7,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits_ctrl_wid,
  output [4:0] io_deq_bits_ctrl_reg_idxw,
  output       io_deq_bits_ctrl_wfd,
  output       io_deq_bits_ctrl_wxd,
  output       io_deq_bits_mask_0,
  output       io_deq_bits_mask_1,
  output       io_deq_bits_mask_2,
  output       io_deq_bits_mask_3,
  output       io_deq_bits_mask_4,
  output       io_deq_bits_mask_5,
  output       io_deq_bits_mask_6,
  output       io_deq_bits_mask_7
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_ctrl_wid [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_ctrl_reg_idxw [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_reg_idxw_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wfd [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_wfd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_wfd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wxd [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_wxd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_ctrl_wxd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_0 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_1 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_2 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_3 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_4 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_5 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_6 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_7 [0:4]; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = enq_ptr_value == 3'h4; // @[Counter.scala 74:24]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  wire  _GEN_53 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_53 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  wrap_1 = deq_ptr_value == 3'h4; // @[Counter.scala 74:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_ctrl_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wid_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_wid_io_deq_bits_MPORT_data = ram_ctrl_wid[ram_ctrl_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_ctrl_wid_io_deq_bits_MPORT_data = ram_ctrl_wid_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_1[1:0] :
    ram_ctrl_wid[ram_ctrl_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_wid_MPORT_data = io_enq_bits_ctrl_wid;
  assign ram_ctrl_wid_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_wid_MPORT_mask = 1'h1;
  assign ram_ctrl_wid_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_data = ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_data = ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_3[4:0] :
    ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_reg_idxw_MPORT_data = io_enq_bits_ctrl_reg_idxw;
  assign ram_ctrl_reg_idxw_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_reg_idxw_MPORT_mask = 1'h1;
  assign ram_ctrl_reg_idxw_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_wfd_io_deq_bits_MPORT_data = ram_ctrl_wfd[ram_ctrl_wfd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_ctrl_wfd_io_deq_bits_MPORT_data = ram_ctrl_wfd_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_5[0:0] :
    ram_ctrl_wfd[ram_ctrl_wfd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_wfd_MPORT_data = io_enq_bits_ctrl_wfd;
  assign ram_ctrl_wfd_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_wfd_MPORT_mask = 1'h1;
  assign ram_ctrl_wfd_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_wxd_io_deq_bits_MPORT_data = ram_ctrl_wxd[ram_ctrl_wxd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_ctrl_wxd_io_deq_bits_MPORT_data = ram_ctrl_wxd_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_7[0:0] :
    ram_ctrl_wxd[ram_ctrl_wxd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ctrl_wxd_MPORT_data = io_enq_bits_ctrl_wxd;
  assign ram_ctrl_wxd_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_wxd_MPORT_mask = 1'h1;
  assign ram_ctrl_wxd_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_0_io_deq_bits_MPORT_data = ram_mask_0[ram_mask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_0_io_deq_bits_MPORT_data = ram_mask_0_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_9[0:0] :
    ram_mask_0[ram_mask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_0_MPORT_data = io_enq_bits_mask_0;
  assign ram_mask_0_MPORT_addr = enq_ptr_value;
  assign ram_mask_0_MPORT_mask = 1'h1;
  assign ram_mask_0_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_1_io_deq_bits_MPORT_data = ram_mask_1[ram_mask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_1_io_deq_bits_MPORT_data = ram_mask_1_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_11[0:0] :
    ram_mask_1[ram_mask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_1_MPORT_data = io_enq_bits_mask_1;
  assign ram_mask_1_MPORT_addr = enq_ptr_value;
  assign ram_mask_1_MPORT_mask = 1'h1;
  assign ram_mask_1_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_2_io_deq_bits_MPORT_data = ram_mask_2[ram_mask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_2_io_deq_bits_MPORT_data = ram_mask_2_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_13[0:0] :
    ram_mask_2[ram_mask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_2_MPORT_data = io_enq_bits_mask_2;
  assign ram_mask_2_MPORT_addr = enq_ptr_value;
  assign ram_mask_2_MPORT_mask = 1'h1;
  assign ram_mask_2_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_3_io_deq_bits_MPORT_data = ram_mask_3[ram_mask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_3_io_deq_bits_MPORT_data = ram_mask_3_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_15[0:0] :
    ram_mask_3[ram_mask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_3_MPORT_data = io_enq_bits_mask_3;
  assign ram_mask_3_MPORT_addr = enq_ptr_value;
  assign ram_mask_3_MPORT_mask = 1'h1;
  assign ram_mask_3_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_4_io_deq_bits_MPORT_data = ram_mask_4[ram_mask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_4_io_deq_bits_MPORT_data = ram_mask_4_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_17[0:0] :
    ram_mask_4[ram_mask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_4_MPORT_data = io_enq_bits_mask_4;
  assign ram_mask_4_MPORT_addr = enq_ptr_value;
  assign ram_mask_4_MPORT_mask = 1'h1;
  assign ram_mask_4_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_5_io_deq_bits_MPORT_data = ram_mask_5[ram_mask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_5_io_deq_bits_MPORT_data = ram_mask_5_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_19[0:0] :
    ram_mask_5[ram_mask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_5_MPORT_data = io_enq_bits_mask_5;
  assign ram_mask_5_MPORT_addr = enq_ptr_value;
  assign ram_mask_5_MPORT_mask = 1'h1;
  assign ram_mask_5_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_6_io_deq_bits_MPORT_data = ram_mask_6[ram_mask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_6_io_deq_bits_MPORT_data = ram_mask_6_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_21[0:0] :
    ram_mask_6[ram_mask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_6_MPORT_data = io_enq_bits_mask_6;
  assign ram_mask_6_MPORT_addr = enq_ptr_value;
  assign ram_mask_6_MPORT_mask = 1'h1;
  assign ram_mask_6_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign ram_mask_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_7_io_deq_bits_MPORT_data = ram_mask_7[ram_mask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_mask_7_io_deq_bits_MPORT_data = ram_mask_7_io_deq_bits_MPORT_addr >= 3'h5 ? _RAND_23[0:0] :
    ram_mask_7[ram_mask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mask_7_MPORT_data = io_enq_bits_mask_7;
  assign ram_mask_7_MPORT_addr = enq_ptr_value;
  assign ram_mask_7_MPORT_mask = 1'h1;
  assign ram_mask_7_MPORT_en = empty ? _GEN_53 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_ctrl_wid = empty ? io_enq_bits_ctrl_wid : ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_ctrl_reg_idxw = empty ? io_enq_bits_ctrl_reg_idxw : ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_ctrl_wfd = empty ? io_enq_bits_ctrl_wfd : ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_ctrl_wxd = empty ? io_enq_bits_ctrl_wxd : ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_0 = empty ? io_enq_bits_mask_0 : ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_1 = empty ? io_enq_bits_mask_1 : ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_2 = empty ? io_enq_bits_mask_2 : ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_3 = empty ? io_enq_bits_mask_3 : ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_4 = empty ? io_enq_bits_mask_4 : ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_5 = empty ? io_enq_bits_mask_5 : ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_6 = empty ? io_enq_bits_mask_6 : ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_7 = empty ? io_enq_bits_mask_7 : ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_ctrl_wid_MPORT_en & ram_ctrl_wid_MPORT_mask) begin
      ram_ctrl_wid[ram_ctrl_wid_MPORT_addr] <= ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_reg_idxw_MPORT_en & ram_ctrl_reg_idxw_MPORT_mask) begin
      ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_MPORT_addr] <= ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wfd_MPORT_en & ram_ctrl_wfd_MPORT_mask) begin
      ram_ctrl_wfd[ram_ctrl_wfd_MPORT_addr] <= ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wxd_MPORT_en & ram_ctrl_wxd_MPORT_mask) begin
      ram_ctrl_wxd[ram_ctrl_wxd_MPORT_addr] <= ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_0_MPORT_en & ram_mask_0_MPORT_mask) begin
      ram_mask_0[ram_mask_0_MPORT_addr] <= ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_1_MPORT_en & ram_mask_1_MPORT_mask) begin
      ram_mask_1[ram_mask_1_MPORT_addr] <= ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_2_MPORT_en & ram_mask_2_MPORT_mask) begin
      ram_mask_2[ram_mask_2_MPORT_addr] <= ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_3_MPORT_en & ram_mask_3_MPORT_mask) begin
      ram_mask_3[ram_mask_3_MPORT_addr] <= ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_4_MPORT_en & ram_mask_4_MPORT_mask) begin
      ram_mask_4[ram_mask_4_MPORT_addr] <= ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_5_MPORT_en & ram_mask_5_MPORT_mask) begin
      ram_mask_5[ram_mask_5_MPORT_addr] <= ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_6_MPORT_en & ram_mask_6_MPORT_mask) begin
      ram_mask_6[ram_mask_6_MPORT_addr] <= ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_7_MPORT_en & ram_mask_7_MPORT_mask) begin
      ram_mask_7[ram_mask_7_MPORT_addr] <= ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      if (wrap) begin // @[Counter.scala 88:20]
        enq_ptr_value <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      if (wrap_1) begin // @[Counter.scala 88:20]
        deq_ptr_value <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
  _RAND_17 = {1{`RANDOM}};
  _RAND_19 = {1{`RANDOM}};
  _RAND_21 = {1{`RANDOM}};
  _RAND_23 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_ctrl_wid[initvar] = _RAND_0[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_ctrl_reg_idxw[initvar] = _RAND_2[4:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_ctrl_wfd[initvar] = _RAND_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_ctrl_wxd[initvar] = _RAND_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_0[initvar] = _RAND_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_1[initvar] = _RAND_10[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_2[initvar] = _RAND_12[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_3[initvar] = _RAND_14[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_4[initvar] = _RAND_16[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_5[initvar] = _RAND_18[0:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_6[initvar] = _RAND_20[0:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    ram_mask_7[initvar] = _RAND_22[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  enq_ptr_value = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  deq_ptr_value = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  maybe_full = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_40(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits_ctrl_wid,
  input  [4:0] io_enq_bits_ctrl_reg_idxw,
  input        io_enq_bits_ctrl_wfd,
  input        io_enq_bits_ctrl_wxd,
  input        io_enq_bits_mask_0,
  input        io_enq_bits_mask_1,
  input        io_enq_bits_mask_2,
  input        io_enq_bits_mask_3,
  input        io_enq_bits_mask_4,
  input        io_enq_bits_mask_5,
  input        io_enq_bits_mask_6,
  input        io_enq_bits_mask_7,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits_ctrl_wid,
  output [4:0] io_deq_bits_ctrl_reg_idxw,
  output       io_deq_bits_ctrl_wfd,
  output       io_deq_bits_ctrl_wxd,
  output       io_deq_bits_mask_0,
  output       io_deq_bits_mask_1,
  output       io_deq_bits_mask_2,
  output       io_deq_bits_mask_3,
  output       io_deq_bits_mask_4,
  output       io_deq_bits_mask_5,
  output       io_deq_bits_mask_6,
  output       io_deq_bits_mask_7
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_ctrl_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_ctrl_reg_idxw [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wfd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wxd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_48 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_48 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_ctrl_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wid_io_deq_bits_MPORT_data = ram_ctrl_wid[ram_ctrl_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wid_MPORT_data = io_enq_bits_ctrl_wid;
  assign ram_ctrl_wid_MPORT_addr = 1'h0;
  assign ram_ctrl_wid_MPORT_mask = 1'h1;
  assign ram_ctrl_wid_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_data = ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_reg_idxw_MPORT_data = io_enq_bits_ctrl_reg_idxw;
  assign ram_ctrl_reg_idxw_MPORT_addr = 1'h0;
  assign ram_ctrl_reg_idxw_MPORT_mask = 1'h1;
  assign ram_ctrl_reg_idxw_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_data = ram_ctrl_wfd[ram_ctrl_wfd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wfd_MPORT_data = io_enq_bits_ctrl_wfd;
  assign ram_ctrl_wfd_MPORT_addr = 1'h0;
  assign ram_ctrl_wfd_MPORT_mask = 1'h1;
  assign ram_ctrl_wfd_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_data = ram_ctrl_wxd[ram_ctrl_wxd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wxd_MPORT_data = io_enq_bits_ctrl_wxd;
  assign ram_ctrl_wxd_MPORT_addr = 1'h0;
  assign ram_ctrl_wxd_MPORT_mask = 1'h1;
  assign ram_ctrl_wxd_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_0_io_deq_bits_MPORT_data = ram_mask_0[ram_mask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_0_MPORT_data = io_enq_bits_mask_0;
  assign ram_mask_0_MPORT_addr = 1'h0;
  assign ram_mask_0_MPORT_mask = 1'h1;
  assign ram_mask_0_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_1_io_deq_bits_MPORT_data = ram_mask_1[ram_mask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_1_MPORT_data = io_enq_bits_mask_1;
  assign ram_mask_1_MPORT_addr = 1'h0;
  assign ram_mask_1_MPORT_mask = 1'h1;
  assign ram_mask_1_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_2_io_deq_bits_MPORT_data = ram_mask_2[ram_mask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_2_MPORT_data = io_enq_bits_mask_2;
  assign ram_mask_2_MPORT_addr = 1'h0;
  assign ram_mask_2_MPORT_mask = 1'h1;
  assign ram_mask_2_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_3_io_deq_bits_MPORT_data = ram_mask_3[ram_mask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_3_MPORT_data = io_enq_bits_mask_3;
  assign ram_mask_3_MPORT_addr = 1'h0;
  assign ram_mask_3_MPORT_mask = 1'h1;
  assign ram_mask_3_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_4_io_deq_bits_MPORT_data = ram_mask_4[ram_mask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_4_MPORT_data = io_enq_bits_mask_4;
  assign ram_mask_4_MPORT_addr = 1'h0;
  assign ram_mask_4_MPORT_mask = 1'h1;
  assign ram_mask_4_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_5_io_deq_bits_MPORT_data = ram_mask_5[ram_mask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_5_MPORT_data = io_enq_bits_mask_5;
  assign ram_mask_5_MPORT_addr = 1'h0;
  assign ram_mask_5_MPORT_mask = 1'h1;
  assign ram_mask_5_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_6_io_deq_bits_MPORT_data = ram_mask_6[ram_mask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_6_MPORT_data = io_enq_bits_mask_6;
  assign ram_mask_6_MPORT_addr = 1'h0;
  assign ram_mask_6_MPORT_mask = 1'h1;
  assign ram_mask_6_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign ram_mask_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_7_io_deq_bits_MPORT_data = ram_mask_7[ram_mask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_7_MPORT_data = io_enq_bits_mask_7;
  assign ram_mask_7_MPORT_addr = 1'h0;
  assign ram_mask_7_MPORT_mask = 1'h1;
  assign ram_mask_7_MPORT_en = empty ? _GEN_48 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_ctrl_wid = empty ? io_enq_bits_ctrl_wid : ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_ctrl_reg_idxw = empty ? io_enq_bits_ctrl_reg_idxw : ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_ctrl_wfd = empty ? io_enq_bits_ctrl_wfd : ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_ctrl_wxd = empty ? io_enq_bits_ctrl_wxd : ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_0 = empty ? io_enq_bits_mask_0 : ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_1 = empty ? io_enq_bits_mask_1 : ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_2 = empty ? io_enq_bits_mask_2 : ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_3 = empty ? io_enq_bits_mask_3 : ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_4 = empty ? io_enq_bits_mask_4 : ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_5 = empty ? io_enq_bits_mask_5 : ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_6 = empty ? io_enq_bits_mask_6 : ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_7 = empty ? io_enq_bits_mask_7 : ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_ctrl_wid_MPORT_en & ram_ctrl_wid_MPORT_mask) begin
      ram_ctrl_wid[ram_ctrl_wid_MPORT_addr] <= ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_reg_idxw_MPORT_en & ram_ctrl_reg_idxw_MPORT_mask) begin
      ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_MPORT_addr] <= ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wfd_MPORT_en & ram_ctrl_wfd_MPORT_mask) begin
      ram_ctrl_wfd[ram_ctrl_wfd_MPORT_addr] <= ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wxd_MPORT_en & ram_ctrl_wxd_MPORT_mask) begin
      ram_ctrl_wxd[ram_ctrl_wxd_MPORT_addr] <= ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_0_MPORT_en & ram_mask_0_MPORT_mask) begin
      ram_mask_0[ram_mask_0_MPORT_addr] <= ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_1_MPORT_en & ram_mask_1_MPORT_mask) begin
      ram_mask_1[ram_mask_1_MPORT_addr] <= ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_2_MPORT_en & ram_mask_2_MPORT_mask) begin
      ram_mask_2[ram_mask_2_MPORT_addr] <= ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_3_MPORT_en & ram_mask_3_MPORT_mask) begin
      ram_mask_3[ram_mask_3_MPORT_addr] <= ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_4_MPORT_en & ram_mask_4_MPORT_mask) begin
      ram_mask_4[ram_mask_4_MPORT_addr] <= ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_5_MPORT_en & ram_mask_5_MPORT_mask) begin
      ram_mask_5[ram_mask_5_MPORT_addr] <= ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_6_MPORT_en & ram_mask_6_MPORT_mask) begin
      ram_mask_6[ram_mask_6_MPORT_addr] <= ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_7_MPORT_en & ram_mask_7_MPORT_mask) begin
      ram_mask_7[ram_mask_7_MPORT_addr] <= ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wid[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_reg_idxw[initvar] = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wfd[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wxd[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_0[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_1[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_2[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_3[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_4[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_5[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_6[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_7[initvar] = _RAND_11[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  maybe_full = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPUexe(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_in1_0,
  input  [31:0] io_in_bits_in1_1,
  input  [31:0] io_in_bits_in1_2,
  input  [31:0] io_in_bits_in1_3,
  input  [31:0] io_in_bits_in1_4,
  input  [31:0] io_in_bits_in1_5,
  input  [31:0] io_in_bits_in1_6,
  input  [31:0] io_in_bits_in1_7,
  input  [31:0] io_in_bits_in2_0,
  input  [31:0] io_in_bits_in2_1,
  input  [31:0] io_in_bits_in2_2,
  input  [31:0] io_in_bits_in2_3,
  input  [31:0] io_in_bits_in2_4,
  input  [31:0] io_in_bits_in2_5,
  input  [31:0] io_in_bits_in2_6,
  input  [31:0] io_in_bits_in2_7,
  input  [31:0] io_in_bits_in3_0,
  input  [31:0] io_in_bits_in3_1,
  input  [31:0] io_in_bits_in3_2,
  input  [31:0] io_in_bits_in3_3,
  input  [31:0] io_in_bits_in3_4,
  input  [31:0] io_in_bits_in3_5,
  input  [31:0] io_in_bits_in3_6,
  input  [31:0] io_in_bits_in3_7,
  input         io_in_bits_mask_0,
  input         io_in_bits_mask_1,
  input         io_in_bits_mask_2,
  input         io_in_bits_mask_3,
  input         io_in_bits_mask_4,
  input         io_in_bits_mask_5,
  input         io_in_bits_mask_6,
  input         io_in_bits_mask_7,
  input  [1:0]  io_in_bits_ctrl_wid,
  input         io_in_bits_ctrl_reverse,
  input  [5:0]  io_in_bits_ctrl_alu_fn,
  input  [4:0]  io_in_bits_ctrl_reg_idxw,
  input         io_in_bits_ctrl_wfd,
  input         io_in_bits_ctrl_wxd,
  input  [2:0]  io_rm,
  input         io_out_x_ready,
  output        io_out_x_valid,
  output [31:0] io_out_x_bits_wb_wxd_rd,
  output        io_out_x_bits_wxd,
  output [4:0]  io_out_x_bits_reg_idxw,
  output [1:0]  io_out_x_bits_warp_id,
  input         io_out_v_ready,
  output        io_out_v_valid,
  output [31:0] io_out_v_bits_wb_wfd_rd_0,
  output [31:0] io_out_v_bits_wb_wfd_rd_1,
  output [31:0] io_out_v_bits_wb_wfd_rd_2,
  output [31:0] io_out_v_bits_wb_wfd_rd_3,
  output [31:0] io_out_v_bits_wb_wfd_rd_4,
  output [31:0] io_out_v_bits_wb_wfd_rd_5,
  output [31:0] io_out_v_bits_wb_wfd_rd_6,
  output [31:0] io_out_v_bits_wb_wfd_rd_7,
  output        io_out_v_bits_wfd_mask_0,
  output        io_out_v_bits_wfd_mask_1,
  output        io_out_v_bits_wfd_mask_2,
  output        io_out_v_bits_wfd_mask_3,
  output        io_out_v_bits_wfd_mask_4,
  output        io_out_v_bits_wfd_mask_5,
  output        io_out_v_bits_wfd_mask_6,
  output        io_out_v_bits_wfd_mask_7,
  output        io_out_v_bits_wfd,
  output [4:0]  io_out_v_bits_reg_idxw,
  output [1:0]  io_out_v_bits_warp_id
);
  wire  ScalarFPU_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_1_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_1_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_1_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_1_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_1_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_1_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_1_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_1_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_1_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_1_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_1_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_1_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_1_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_2_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_2_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_2_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_2_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_2_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_2_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_2_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_2_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_2_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_2_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_2_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_2_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_2_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_3_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_3_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_3_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_3_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_3_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_3_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_3_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_3_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_3_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_3_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_3_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_3_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_3_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_4_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_4_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_4_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_4_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_4_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_4_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_4_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_4_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_4_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_4_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_4_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_4_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_4_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_5_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_5_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_5_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_5_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_5_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_5_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_5_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_5_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_5_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_5_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_5_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_5_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_5_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_6_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_6_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_6_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_6_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_6_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_6_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_6_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_6_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_6_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_6_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_6_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_6_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_6_io_select; // @[execution.scala 114:47]
  wire  ScalarFPU_7_clock; // @[execution.scala 114:47]
  wire  ScalarFPU_7_reset; // @[execution.scala 114:47]
  wire  ScalarFPU_7_io_in_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_7_io_in_valid; // @[execution.scala 114:47]
  wire [5:0] ScalarFPU_7_io_in_bits_fpuop; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_7_io_in_bits_a; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_7_io_in_bits_b; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_7_io_in_bits_c; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_7_io_in_bits_rm; // @[execution.scala 114:47]
  wire  ScalarFPU_7_io_out_ready; // @[execution.scala 114:47]
  wire  ScalarFPU_7_io_out_valid; // @[execution.scala 114:47]
  wire [31:0] ScalarFPU_7_io_out_bits_result; // @[execution.scala 114:47]
  wire [2:0] ScalarFPU_7_io_select; // @[execution.scala 114:47]
  wire  result_x_clock; // @[execution.scala 115:22]
  wire  result_x_reset; // @[execution.scala 115:22]
  wire  result_x_io_enq_ready; // @[execution.scala 115:22]
  wire  result_x_io_enq_valid; // @[execution.scala 115:22]
  wire [31:0] result_x_io_enq_bits_wb_wxd_rd; // @[execution.scala 115:22]
  wire  result_x_io_enq_bits_wxd; // @[execution.scala 115:22]
  wire [4:0] result_x_io_enq_bits_reg_idxw; // @[execution.scala 115:22]
  wire [1:0] result_x_io_enq_bits_warp_id; // @[execution.scala 115:22]
  wire  result_x_io_deq_ready; // @[execution.scala 115:22]
  wire  result_x_io_deq_valid; // @[execution.scala 115:22]
  wire [31:0] result_x_io_deq_bits_wb_wxd_rd; // @[execution.scala 115:22]
  wire  result_x_io_deq_bits_wxd; // @[execution.scala 115:22]
  wire [4:0] result_x_io_deq_bits_reg_idxw; // @[execution.scala 115:22]
  wire [1:0] result_x_io_deq_bits_warp_id; // @[execution.scala 115:22]
  wire  result_v_clock; // @[execution.scala 116:22]
  wire  result_v_reset; // @[execution.scala 116:22]
  wire  result_v_io_enq_ready; // @[execution.scala 116:22]
  wire  result_v_io_enq_valid; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_0; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_1; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_2; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_3; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_4; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_5; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_6; // @[execution.scala 116:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_7; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_0; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_1; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_2; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_3; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_4; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_5; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_6; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd_mask_7; // @[execution.scala 116:22]
  wire  result_v_io_enq_bits_wfd; // @[execution.scala 116:22]
  wire [4:0] result_v_io_enq_bits_reg_idxw; // @[execution.scala 116:22]
  wire [1:0] result_v_io_enq_bits_warp_id; // @[execution.scala 116:22]
  wire  result_v_io_deq_ready; // @[execution.scala 116:22]
  wire  result_v_io_deq_valid; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_0; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_1; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_2; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_3; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_4; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_5; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_6; // @[execution.scala 116:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_7; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_0; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_1; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_2; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_3; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_4; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_5; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_6; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd_mask_7; // @[execution.scala 116:22]
  wire  result_v_io_deq_bits_wfd; // @[execution.scala 116:22]
  wire [4:0] result_v_io_deq_bits_reg_idxw; // @[execution.scala 116:22]
  wire [1:0] result_v_io_deq_bits_warp_id; // @[execution.scala 116:22]
  wire  ctrl_fma_clock; // @[execution.scala 138:22]
  wire  ctrl_fma_reset; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_ready; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_valid; // @[execution.scala 138:22]
  wire [1:0] ctrl_fma_io_enq_bits_ctrl_wid; // @[execution.scala 138:22]
  wire [4:0] ctrl_fma_io_enq_bits_ctrl_reg_idxw; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_ctrl_wfd; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_ctrl_wxd; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_0; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_1; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_2; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_3; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_4; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_5; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_6; // @[execution.scala 138:22]
  wire  ctrl_fma_io_enq_bits_mask_7; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_ready; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_valid; // @[execution.scala 138:22]
  wire [1:0] ctrl_fma_io_deq_bits_ctrl_wid; // @[execution.scala 138:22]
  wire [4:0] ctrl_fma_io_deq_bits_ctrl_reg_idxw; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_ctrl_wfd; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_ctrl_wxd; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_0; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_1; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_2; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_3; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_4; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_5; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_6; // @[execution.scala 138:22]
  wire  ctrl_fma_io_deq_bits_mask_7; // @[execution.scala 138:22]
  wire  ctrl_else_clock; // @[execution.scala 139:23]
  wire  ctrl_else_reset; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_ready; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_valid; // @[execution.scala 139:23]
  wire [1:0] ctrl_else_io_enq_bits_ctrl_wid; // @[execution.scala 139:23]
  wire [4:0] ctrl_else_io_enq_bits_ctrl_reg_idxw; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_ctrl_wfd; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_ctrl_wxd; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_0; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_1; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_2; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_3; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_4; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_5; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_6; // @[execution.scala 139:23]
  wire  ctrl_else_io_enq_bits_mask_7; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_ready; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_valid; // @[execution.scala 139:23]
  wire [1:0] ctrl_else_io_deq_bits_ctrl_wid; // @[execution.scala 139:23]
  wire [4:0] ctrl_else_io_deq_bits_ctrl_reg_idxw; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_ctrl_wfd; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_ctrl_wxd; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_0; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_1; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_2; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_3; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_4; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_5; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_6; // @[execution.scala 139:23]
  wire  ctrl_else_io_deq_bits_mask_7; // @[execution.scala 139:23]
  wire [31:0] _GEN_0 = io_in_bits_ctrl_reverse ? io_in_bits_in2_0 : io_in_bits_in1_0; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_1 = io_in_bits_ctrl_reverse ? io_in_bits_in1_0 : io_in_bits_in2_0; // @[execution.scala 119:22 126:35 128:24]
  wire [5:0] _fpu_0_in_bits_fpuop_T_1 = io_in_bits_ctrl_alu_fn - 6'ha; // @[execution.scala 131:51]
  wire [5:0] fpu_0_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  wire [31:0] _GEN_6 = io_in_bits_ctrl_reverse ? io_in_bits_in2_1 : io_in_bits_in1_1; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_7 = io_in_bits_ctrl_reverse ? io_in_bits_in1_1 : io_in_bits_in2_1; // @[execution.scala 119:22 126:35 128:24]
  wire [31:0] _GEN_12 = io_in_bits_ctrl_reverse ? io_in_bits_in2_2 : io_in_bits_in1_2; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_13 = io_in_bits_ctrl_reverse ? io_in_bits_in1_2 : io_in_bits_in2_2; // @[execution.scala 119:22 126:35 128:24]
  wire [31:0] _GEN_18 = io_in_bits_ctrl_reverse ? io_in_bits_in2_3 : io_in_bits_in1_3; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_19 = io_in_bits_ctrl_reverse ? io_in_bits_in1_3 : io_in_bits_in2_3; // @[execution.scala 119:22 126:35 128:24]
  wire [31:0] _GEN_24 = io_in_bits_ctrl_reverse ? io_in_bits_in2_4 : io_in_bits_in1_4; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_25 = io_in_bits_ctrl_reverse ? io_in_bits_in1_4 : io_in_bits_in2_4; // @[execution.scala 119:22 126:35 128:24]
  wire [31:0] _GEN_30 = io_in_bits_ctrl_reverse ? io_in_bits_in2_5 : io_in_bits_in1_5; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_31 = io_in_bits_ctrl_reverse ? io_in_bits_in1_5 : io_in_bits_in2_5; // @[execution.scala 119:22 126:35 128:24]
  wire [31:0] _GEN_36 = io_in_bits_ctrl_reverse ? io_in_bits_in2_6 : io_in_bits_in1_6; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_37 = io_in_bits_ctrl_reverse ? io_in_bits_in1_6 : io_in_bits_in2_6; // @[execution.scala 119:22 126:35 128:24]
  wire [31:0] _GEN_42 = io_in_bits_ctrl_reverse ? io_in_bits_in2_7 : io_in_bits_in1_7; // @[execution.scala 118:22 126:35 127:24]
  wire [31:0] _GEN_43 = io_in_bits_ctrl_reverse ? io_in_bits_in1_7 : io_in_bits_in2_7; // @[execution.scala 119:22 126:35 128:24]
  wire  fpu_0_in_ready = ScalarFPU_io_in_ready; // @[execution.scala 114:{18,18}]
  wire  _ctrl_fma_io_enq_valid_T = fpu_0_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  wire [2:0] fpu_0_select = ScalarFPU_io_select; // @[execution.scala 114:{18,18}]
  wire  _ctrl_T = fpu_0_select == 3'h0; // @[execution.scala 148:29]
  wire  ctrl_ctrl_wxd = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_wxd : ctrl_else_io_deq_bits_ctrl_wxd; // @[execution.scala 148:15]
  wire  fpu_0_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  wire  fpu_0_out_valid = ScalarFPU_io_out_valid; // @[execution.scala 114:{18,18}]
  wire  _ctrl_fma_io_deq_ready_T = fpu_0_out_ready & fpu_0_out_valid; // @[Decoupled.scala 50:35]
  wire  ctrl_ctrl_wfd = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_wfd : ctrl_else_io_deq_bits_ctrl_wfd; // @[execution.scala 148:15]
  ScalarFPU ScalarFPU ( // @[execution.scala 114:47]
    .clock(ScalarFPU_clock),
    .reset(ScalarFPU_reset),
    .io_in_ready(ScalarFPU_io_in_ready),
    .io_in_valid(ScalarFPU_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_io_in_bits_rm),
    .io_out_ready(ScalarFPU_io_out_ready),
    .io_out_valid(ScalarFPU_io_out_valid),
    .io_out_bits_result(ScalarFPU_io_out_bits_result),
    .io_select(ScalarFPU_io_select)
  );
  ScalarFPU ScalarFPU_1 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_1_clock),
    .reset(ScalarFPU_1_reset),
    .io_in_ready(ScalarFPU_1_io_in_ready),
    .io_in_valid(ScalarFPU_1_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_1_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_1_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_1_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_1_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_1_io_in_bits_rm),
    .io_out_ready(ScalarFPU_1_io_out_ready),
    .io_out_valid(ScalarFPU_1_io_out_valid),
    .io_out_bits_result(ScalarFPU_1_io_out_bits_result),
    .io_select(ScalarFPU_1_io_select)
  );
  ScalarFPU ScalarFPU_2 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_2_clock),
    .reset(ScalarFPU_2_reset),
    .io_in_ready(ScalarFPU_2_io_in_ready),
    .io_in_valid(ScalarFPU_2_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_2_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_2_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_2_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_2_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_2_io_in_bits_rm),
    .io_out_ready(ScalarFPU_2_io_out_ready),
    .io_out_valid(ScalarFPU_2_io_out_valid),
    .io_out_bits_result(ScalarFPU_2_io_out_bits_result),
    .io_select(ScalarFPU_2_io_select)
  );
  ScalarFPU ScalarFPU_3 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_3_clock),
    .reset(ScalarFPU_3_reset),
    .io_in_ready(ScalarFPU_3_io_in_ready),
    .io_in_valid(ScalarFPU_3_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_3_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_3_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_3_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_3_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_3_io_in_bits_rm),
    .io_out_ready(ScalarFPU_3_io_out_ready),
    .io_out_valid(ScalarFPU_3_io_out_valid),
    .io_out_bits_result(ScalarFPU_3_io_out_bits_result),
    .io_select(ScalarFPU_3_io_select)
  );
  ScalarFPU ScalarFPU_4 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_4_clock),
    .reset(ScalarFPU_4_reset),
    .io_in_ready(ScalarFPU_4_io_in_ready),
    .io_in_valid(ScalarFPU_4_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_4_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_4_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_4_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_4_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_4_io_in_bits_rm),
    .io_out_ready(ScalarFPU_4_io_out_ready),
    .io_out_valid(ScalarFPU_4_io_out_valid),
    .io_out_bits_result(ScalarFPU_4_io_out_bits_result),
    .io_select(ScalarFPU_4_io_select)
  );
  ScalarFPU ScalarFPU_5 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_5_clock),
    .reset(ScalarFPU_5_reset),
    .io_in_ready(ScalarFPU_5_io_in_ready),
    .io_in_valid(ScalarFPU_5_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_5_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_5_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_5_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_5_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_5_io_in_bits_rm),
    .io_out_ready(ScalarFPU_5_io_out_ready),
    .io_out_valid(ScalarFPU_5_io_out_valid),
    .io_out_bits_result(ScalarFPU_5_io_out_bits_result),
    .io_select(ScalarFPU_5_io_select)
  );
  ScalarFPU ScalarFPU_6 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_6_clock),
    .reset(ScalarFPU_6_reset),
    .io_in_ready(ScalarFPU_6_io_in_ready),
    .io_in_valid(ScalarFPU_6_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_6_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_6_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_6_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_6_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_6_io_in_bits_rm),
    .io_out_ready(ScalarFPU_6_io_out_ready),
    .io_out_valid(ScalarFPU_6_io_out_valid),
    .io_out_bits_result(ScalarFPU_6_io_out_bits_result),
    .io_select(ScalarFPU_6_io_select)
  );
  ScalarFPU ScalarFPU_7 ( // @[execution.scala 114:47]
    .clock(ScalarFPU_7_clock),
    .reset(ScalarFPU_7_reset),
    .io_in_ready(ScalarFPU_7_io_in_ready),
    .io_in_valid(ScalarFPU_7_io_in_valid),
    .io_in_bits_fpuop(ScalarFPU_7_io_in_bits_fpuop),
    .io_in_bits_a(ScalarFPU_7_io_in_bits_a),
    .io_in_bits_b(ScalarFPU_7_io_in_bits_b),
    .io_in_bits_c(ScalarFPU_7_io_in_bits_c),
    .io_in_bits_rm(ScalarFPU_7_io_in_bits_rm),
    .io_out_ready(ScalarFPU_7_io_out_ready),
    .io_out_valid(ScalarFPU_7_io_out_valid),
    .io_out_bits_result(ScalarFPU_7_io_out_bits_result),
    .io_select(ScalarFPU_7_io_select)
  );
  Queue_1 result_x ( // @[execution.scala 115:22]
    .clock(result_x_clock),
    .reset(result_x_reset),
    .io_enq_ready(result_x_io_enq_ready),
    .io_enq_valid(result_x_io_enq_valid),
    .io_enq_bits_wb_wxd_rd(result_x_io_enq_bits_wb_wxd_rd),
    .io_enq_bits_wxd(result_x_io_enq_bits_wxd),
    .io_enq_bits_reg_idxw(result_x_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_x_io_enq_bits_warp_id),
    .io_deq_ready(result_x_io_deq_ready),
    .io_deq_valid(result_x_io_deq_valid),
    .io_deq_bits_wb_wxd_rd(result_x_io_deq_bits_wb_wxd_rd),
    .io_deq_bits_wxd(result_x_io_deq_bits_wxd),
    .io_deq_bits_reg_idxw(result_x_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_x_io_deq_bits_warp_id)
  );
  Queue_3 result_v ( // @[execution.scala 116:22]
    .clock(result_v_clock),
    .reset(result_v_reset),
    .io_enq_ready(result_v_io_enq_ready),
    .io_enq_valid(result_v_io_enq_valid),
    .io_enq_bits_wb_wfd_rd_0(result_v_io_enq_bits_wb_wfd_rd_0),
    .io_enq_bits_wb_wfd_rd_1(result_v_io_enq_bits_wb_wfd_rd_1),
    .io_enq_bits_wb_wfd_rd_2(result_v_io_enq_bits_wb_wfd_rd_2),
    .io_enq_bits_wb_wfd_rd_3(result_v_io_enq_bits_wb_wfd_rd_3),
    .io_enq_bits_wb_wfd_rd_4(result_v_io_enq_bits_wb_wfd_rd_4),
    .io_enq_bits_wb_wfd_rd_5(result_v_io_enq_bits_wb_wfd_rd_5),
    .io_enq_bits_wb_wfd_rd_6(result_v_io_enq_bits_wb_wfd_rd_6),
    .io_enq_bits_wb_wfd_rd_7(result_v_io_enq_bits_wb_wfd_rd_7),
    .io_enq_bits_wfd_mask_0(result_v_io_enq_bits_wfd_mask_0),
    .io_enq_bits_wfd_mask_1(result_v_io_enq_bits_wfd_mask_1),
    .io_enq_bits_wfd_mask_2(result_v_io_enq_bits_wfd_mask_2),
    .io_enq_bits_wfd_mask_3(result_v_io_enq_bits_wfd_mask_3),
    .io_enq_bits_wfd_mask_4(result_v_io_enq_bits_wfd_mask_4),
    .io_enq_bits_wfd_mask_5(result_v_io_enq_bits_wfd_mask_5),
    .io_enq_bits_wfd_mask_6(result_v_io_enq_bits_wfd_mask_6),
    .io_enq_bits_wfd_mask_7(result_v_io_enq_bits_wfd_mask_7),
    .io_enq_bits_wfd(result_v_io_enq_bits_wfd),
    .io_enq_bits_reg_idxw(result_v_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_v_io_enq_bits_warp_id),
    .io_deq_ready(result_v_io_deq_ready),
    .io_deq_valid(result_v_io_deq_valid),
    .io_deq_bits_wb_wfd_rd_0(result_v_io_deq_bits_wb_wfd_rd_0),
    .io_deq_bits_wb_wfd_rd_1(result_v_io_deq_bits_wb_wfd_rd_1),
    .io_deq_bits_wb_wfd_rd_2(result_v_io_deq_bits_wb_wfd_rd_2),
    .io_deq_bits_wb_wfd_rd_3(result_v_io_deq_bits_wb_wfd_rd_3),
    .io_deq_bits_wb_wfd_rd_4(result_v_io_deq_bits_wb_wfd_rd_4),
    .io_deq_bits_wb_wfd_rd_5(result_v_io_deq_bits_wb_wfd_rd_5),
    .io_deq_bits_wb_wfd_rd_6(result_v_io_deq_bits_wb_wfd_rd_6),
    .io_deq_bits_wb_wfd_rd_7(result_v_io_deq_bits_wb_wfd_rd_7),
    .io_deq_bits_wfd_mask_0(result_v_io_deq_bits_wfd_mask_0),
    .io_deq_bits_wfd_mask_1(result_v_io_deq_bits_wfd_mask_1),
    .io_deq_bits_wfd_mask_2(result_v_io_deq_bits_wfd_mask_2),
    .io_deq_bits_wfd_mask_3(result_v_io_deq_bits_wfd_mask_3),
    .io_deq_bits_wfd_mask_4(result_v_io_deq_bits_wfd_mask_4),
    .io_deq_bits_wfd_mask_5(result_v_io_deq_bits_wfd_mask_5),
    .io_deq_bits_wfd_mask_6(result_v_io_deq_bits_wfd_mask_6),
    .io_deq_bits_wfd_mask_7(result_v_io_deq_bits_wfd_mask_7),
    .io_deq_bits_wfd(result_v_io_deq_bits_wfd),
    .io_deq_bits_reg_idxw(result_v_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_v_io_deq_bits_warp_id)
  );
  Queue_39 ctrl_fma ( // @[execution.scala 138:22]
    .clock(ctrl_fma_clock),
    .reset(ctrl_fma_reset),
    .io_enq_ready(ctrl_fma_io_enq_ready),
    .io_enq_valid(ctrl_fma_io_enq_valid),
    .io_enq_bits_ctrl_wid(ctrl_fma_io_enq_bits_ctrl_wid),
    .io_enq_bits_ctrl_reg_idxw(ctrl_fma_io_enq_bits_ctrl_reg_idxw),
    .io_enq_bits_ctrl_wfd(ctrl_fma_io_enq_bits_ctrl_wfd),
    .io_enq_bits_ctrl_wxd(ctrl_fma_io_enq_bits_ctrl_wxd),
    .io_enq_bits_mask_0(ctrl_fma_io_enq_bits_mask_0),
    .io_enq_bits_mask_1(ctrl_fma_io_enq_bits_mask_1),
    .io_enq_bits_mask_2(ctrl_fma_io_enq_bits_mask_2),
    .io_enq_bits_mask_3(ctrl_fma_io_enq_bits_mask_3),
    .io_enq_bits_mask_4(ctrl_fma_io_enq_bits_mask_4),
    .io_enq_bits_mask_5(ctrl_fma_io_enq_bits_mask_5),
    .io_enq_bits_mask_6(ctrl_fma_io_enq_bits_mask_6),
    .io_enq_bits_mask_7(ctrl_fma_io_enq_bits_mask_7),
    .io_deq_ready(ctrl_fma_io_deq_ready),
    .io_deq_valid(ctrl_fma_io_deq_valid),
    .io_deq_bits_ctrl_wid(ctrl_fma_io_deq_bits_ctrl_wid),
    .io_deq_bits_ctrl_reg_idxw(ctrl_fma_io_deq_bits_ctrl_reg_idxw),
    .io_deq_bits_ctrl_wfd(ctrl_fma_io_deq_bits_ctrl_wfd),
    .io_deq_bits_ctrl_wxd(ctrl_fma_io_deq_bits_ctrl_wxd),
    .io_deq_bits_mask_0(ctrl_fma_io_deq_bits_mask_0),
    .io_deq_bits_mask_1(ctrl_fma_io_deq_bits_mask_1),
    .io_deq_bits_mask_2(ctrl_fma_io_deq_bits_mask_2),
    .io_deq_bits_mask_3(ctrl_fma_io_deq_bits_mask_3),
    .io_deq_bits_mask_4(ctrl_fma_io_deq_bits_mask_4),
    .io_deq_bits_mask_5(ctrl_fma_io_deq_bits_mask_5),
    .io_deq_bits_mask_6(ctrl_fma_io_deq_bits_mask_6),
    .io_deq_bits_mask_7(ctrl_fma_io_deq_bits_mask_7)
  );
  Queue_40 ctrl_else ( // @[execution.scala 139:23]
    .clock(ctrl_else_clock),
    .reset(ctrl_else_reset),
    .io_enq_ready(ctrl_else_io_enq_ready),
    .io_enq_valid(ctrl_else_io_enq_valid),
    .io_enq_bits_ctrl_wid(ctrl_else_io_enq_bits_ctrl_wid),
    .io_enq_bits_ctrl_reg_idxw(ctrl_else_io_enq_bits_ctrl_reg_idxw),
    .io_enq_bits_ctrl_wfd(ctrl_else_io_enq_bits_ctrl_wfd),
    .io_enq_bits_ctrl_wxd(ctrl_else_io_enq_bits_ctrl_wxd),
    .io_enq_bits_mask_0(ctrl_else_io_enq_bits_mask_0),
    .io_enq_bits_mask_1(ctrl_else_io_enq_bits_mask_1),
    .io_enq_bits_mask_2(ctrl_else_io_enq_bits_mask_2),
    .io_enq_bits_mask_3(ctrl_else_io_enq_bits_mask_3),
    .io_enq_bits_mask_4(ctrl_else_io_enq_bits_mask_4),
    .io_enq_bits_mask_5(ctrl_else_io_enq_bits_mask_5),
    .io_enq_bits_mask_6(ctrl_else_io_enq_bits_mask_6),
    .io_enq_bits_mask_7(ctrl_else_io_enq_bits_mask_7),
    .io_deq_ready(ctrl_else_io_deq_ready),
    .io_deq_valid(ctrl_else_io_deq_valid),
    .io_deq_bits_ctrl_wid(ctrl_else_io_deq_bits_ctrl_wid),
    .io_deq_bits_ctrl_reg_idxw(ctrl_else_io_deq_bits_ctrl_reg_idxw),
    .io_deq_bits_ctrl_wfd(ctrl_else_io_deq_bits_ctrl_wfd),
    .io_deq_bits_ctrl_wxd(ctrl_else_io_deq_bits_ctrl_wxd),
    .io_deq_bits_mask_0(ctrl_else_io_deq_bits_mask_0),
    .io_deq_bits_mask_1(ctrl_else_io_deq_bits_mask_1),
    .io_deq_bits_mask_2(ctrl_else_io_deq_bits_mask_2),
    .io_deq_bits_mask_3(ctrl_else_io_deq_bits_mask_3),
    .io_deq_bits_mask_4(ctrl_else_io_deq_bits_mask_4),
    .io_deq_bits_mask_5(ctrl_else_io_deq_bits_mask_5),
    .io_deq_bits_mask_6(ctrl_else_io_deq_bits_mask_6),
    .io_deq_bits_mask_7(ctrl_else_io_deq_bits_mask_7)
  );
  assign io_in_ready = ScalarFPU_io_in_ready; // @[execution.scala 114:{18,18}]
  assign io_out_x_valid = result_x_io_deq_valid; // @[execution.scala 167:11]
  assign io_out_x_bits_wb_wxd_rd = result_x_io_deq_bits_wb_wxd_rd; // @[execution.scala 167:11]
  assign io_out_x_bits_wxd = result_x_io_deq_bits_wxd; // @[execution.scala 167:11]
  assign io_out_x_bits_reg_idxw = result_x_io_deq_bits_reg_idxw; // @[execution.scala 167:11]
  assign io_out_x_bits_warp_id = result_x_io_deq_bits_warp_id; // @[execution.scala 167:11]
  assign io_out_v_valid = result_v_io_deq_valid; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_0 = result_v_io_deq_bits_wb_wfd_rd_0; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_1 = result_v_io_deq_bits_wb_wfd_rd_1; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_2 = result_v_io_deq_bits_wb_wfd_rd_2; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_3 = result_v_io_deq_bits_wb_wfd_rd_3; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_4 = result_v_io_deq_bits_wb_wfd_rd_4; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_5 = result_v_io_deq_bits_wb_wfd_rd_5; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_6 = result_v_io_deq_bits_wb_wfd_rd_6; // @[execution.scala 166:11]
  assign io_out_v_bits_wb_wfd_rd_7 = result_v_io_deq_bits_wb_wfd_rd_7; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_0 = result_v_io_deq_bits_wfd_mask_0; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_1 = result_v_io_deq_bits_wfd_mask_1; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_2 = result_v_io_deq_bits_wfd_mask_2; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_3 = result_v_io_deq_bits_wfd_mask_3; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_4 = result_v_io_deq_bits_wfd_mask_4; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_5 = result_v_io_deq_bits_wfd_mask_5; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_6 = result_v_io_deq_bits_wfd_mask_6; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd_mask_7 = result_v_io_deq_bits_wfd_mask_7; // @[execution.scala 166:11]
  assign io_out_v_bits_wfd = result_v_io_deq_bits_wfd; // @[execution.scala 166:11]
  assign io_out_v_bits_reg_idxw = result_v_io_deq_bits_reg_idxw; // @[execution.scala 166:11]
  assign io_out_v_bits_warp_id = result_v_io_deq_bits_warp_id; // @[execution.scala 166:11]
  assign ScalarFPU_clock = clock;
  assign ScalarFPU_reset = reset;
  assign ScalarFPU_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_0 : _GEN_0; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_0 : _GEN_1; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_0 : io_in_bits_in3_0; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_1_clock = clock;
  assign ScalarFPU_1_reset = reset;
  assign ScalarFPU_1_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_1_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_1_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_1 : _GEN_6; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_1_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_1 : _GEN_7; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_1_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_1 : io_in_bits_in3_1; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_1_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_1_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_2_clock = clock;
  assign ScalarFPU_2_reset = reset;
  assign ScalarFPU_2_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_2_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_2_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_2 : _GEN_12; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_2_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_2 : _GEN_13; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_2_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_2 : io_in_bits_in3_2; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_2_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_2_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_3_clock = clock;
  assign ScalarFPU_3_reset = reset;
  assign ScalarFPU_3_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_3_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_3_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_3 : _GEN_18; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_3_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_3 : _GEN_19; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_3_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_3 : io_in_bits_in3_3; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_3_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_3_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_4_clock = clock;
  assign ScalarFPU_4_reset = reset;
  assign ScalarFPU_4_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_4_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_4_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_4 : _GEN_24; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_4_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_4 : _GEN_25; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_4_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_4 : io_in_bits_in3_4; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_4_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_4_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_5_clock = clock;
  assign ScalarFPU_5_reset = reset;
  assign ScalarFPU_5_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_5_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_5_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_5 : _GEN_30; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_5_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_5 : _GEN_31; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_5_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_5 : io_in_bits_in3_5; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_5_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_5_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_6_clock = clock;
  assign ScalarFPU_6_reset = reset;
  assign ScalarFPU_6_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_6_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_6_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_6 : _GEN_36; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_6_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_6 : _GEN_37; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_6_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_6 : io_in_bits_in3_6; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_6_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_6_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign ScalarFPU_7_clock = clock;
  assign ScalarFPU_7_reset = reset;
  assign ScalarFPU_7_io_in_valid = io_in_valid; // @[execution.scala 114:18 123:20]
  assign ScalarFPU_7_io_in_bits_fpuop = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? _fpu_0_in_bits_fpuop_T_1 :
    io_in_bits_ctrl_alu_fn; // @[execution.scala 130:160 121:26 131:27]
  assign ScalarFPU_7_io_in_bits_a = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in1_7 : _GEN_42; // @[execution.scala 130:160 132:24]
  assign ScalarFPU_7_io_in_bits_b = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in3_7 : _GEN_43; // @[execution.scala 130:160 133:24]
  assign ScalarFPU_7_io_in_bits_c = io_in_bits_ctrl_alu_fn == 6'he | io_in_bits_ctrl_alu_fn == 6'hf |
    io_in_bits_ctrl_alu_fn == 6'h11 | io_in_bits_ctrl_alu_fn == 6'h10 ? io_in_bits_in2_7 : io_in_bits_in3_7; // @[execution.scala 130:160 120:22 134:24]
  assign ScalarFPU_7_io_in_bits_rm = io_rm; // @[execution.scala 114:18 122:23]
  assign ScalarFPU_7_io_out_ready = ctrl_ctrl_wxd ? result_x_io_enq_ready : result_v_io_enq_ready; // @[execution.scala 150:26]
  assign result_x_clock = clock;
  assign result_x_reset = reset;
  assign result_x_io_enq_valid = fpu_0_out_valid & ctrl_ctrl_wxd; // @[execution.scala 164:42]
  assign result_x_io_enq_bits_wb_wxd_rd = ScalarFPU_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_x_io_enq_bits_wxd = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_wxd :
    ctrl_else_io_deq_bits_ctrl_wxd; // @[execution.scala 148:15]
  assign result_x_io_enq_bits_reg_idxw = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_reg_idxw :
    ctrl_else_io_deq_bits_ctrl_reg_idxw; // @[execution.scala 148:15]
  assign result_x_io_enq_bits_warp_id = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_wid :
    ctrl_else_io_deq_bits_ctrl_wid; // @[execution.scala 148:15]
  assign result_x_io_deq_ready = io_out_x_ready; // @[execution.scala 167:11]
  assign result_v_clock = clock;
  assign result_v_reset = reset;
  assign result_v_io_enq_valid = fpu_0_out_valid & ctrl_ctrl_wfd; // @[execution.scala 163:42]
  assign result_v_io_enq_bits_wb_wfd_rd_0 = ScalarFPU_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_1 = ScalarFPU_1_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_2 = ScalarFPU_2_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_3 = ScalarFPU_3_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_4 = ScalarFPU_4_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_5 = ScalarFPU_5_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_6 = ScalarFPU_6_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wb_wfd_rd_7 = ScalarFPU_7_io_out_bits_result; // @[execution.scala 114:{18,18}]
  assign result_v_io_enq_bits_wfd_mask_0 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_0 :
    ctrl_else_io_deq_bits_mask_0; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_1 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_1 :
    ctrl_else_io_deq_bits_mask_1; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_2 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_2 :
    ctrl_else_io_deq_bits_mask_2; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_3 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_3 :
    ctrl_else_io_deq_bits_mask_3; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_4 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_4 :
    ctrl_else_io_deq_bits_mask_4; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_5 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_5 :
    ctrl_else_io_deq_bits_mask_5; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_6 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_6 :
    ctrl_else_io_deq_bits_mask_6; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd_mask_7 = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_mask_7 :
    ctrl_else_io_deq_bits_mask_7; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_wfd = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_wfd :
    ctrl_else_io_deq_bits_ctrl_wfd; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_reg_idxw = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_reg_idxw :
    ctrl_else_io_deq_bits_ctrl_reg_idxw; // @[execution.scala 148:15]
  assign result_v_io_enq_bits_warp_id = fpu_0_select == 3'h0 ? ctrl_fma_io_deq_bits_ctrl_wid :
    ctrl_else_io_deq_bits_ctrl_wid; // @[execution.scala 148:15]
  assign result_v_io_deq_ready = io_out_v_ready; // @[execution.scala 166:11]
  assign ctrl_fma_clock = clock;
  assign ctrl_fma_reset = reset;
  assign ctrl_fma_io_enq_valid = _ctrl_fma_io_enq_valid_T & fpu_0_in_bits_fpuop[5:3] == 3'h0; // @[execution.scala 142:41]
  assign ctrl_fma_io_enq_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[execution.scala 140:28]
  assign ctrl_fma_io_enq_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[execution.scala 140:28]
  assign ctrl_fma_io_enq_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[execution.scala 140:28]
  assign ctrl_fma_io_enq_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[execution.scala 140:28]
  assign ctrl_fma_io_enq_bits_mask_0 = io_in_bits_mask_0; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_1 = io_in_bits_mask_1; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_2 = io_in_bits_mask_2; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_3 = io_in_bits_mask_3; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_4 = io_in_bits_mask_4; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_5 = io_in_bits_mask_5; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_6 = io_in_bits_mask_6; // @[execution.scala 141:28]
  assign ctrl_fma_io_enq_bits_mask_7 = io_in_bits_mask_7; // @[execution.scala 141:28]
  assign ctrl_fma_io_deq_ready = _ctrl_fma_io_deq_ready_T & _ctrl_T; // @[execution.scala 143:42]
  assign ctrl_else_clock = clock;
  assign ctrl_else_reset = reset;
  assign ctrl_else_io_enq_valid = _ctrl_fma_io_enq_valid_T & fpu_0_in_bits_fpuop[5:3] != 3'h0; // @[execution.scala 146:42]
  assign ctrl_else_io_enq_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[execution.scala 144:29]
  assign ctrl_else_io_enq_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[execution.scala 144:29]
  assign ctrl_else_io_enq_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[execution.scala 144:29]
  assign ctrl_else_io_enq_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[execution.scala 144:29]
  assign ctrl_else_io_enq_bits_mask_0 = io_in_bits_mask_0; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_1 = io_in_bits_mask_1; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_2 = io_in_bits_mask_2; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_3 = io_in_bits_mask_3; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_4 = io_in_bits_mask_4; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_5 = io_in_bits_mask_5; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_6 = io_in_bits_mask_6; // @[execution.scala 145:29]
  assign ctrl_else_io_enq_bits_mask_7 = io_in_bits_mask_7; // @[execution.scala 145:29]
  assign ctrl_else_io_deq_ready = _ctrl_fma_io_deq_ready_T & fpu_0_select != 3'h0; // @[execution.scala 147:43]
endmodule
module Queue_41(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_in1_0,
  input  [31:0] io_enq_bits_in1_1,
  input  [31:0] io_enq_bits_in1_2,
  input  [31:0] io_enq_bits_in1_3,
  input  [31:0] io_enq_bits_in1_4,
  input  [31:0] io_enq_bits_in1_5,
  input  [31:0] io_enq_bits_in1_6,
  input  [31:0] io_enq_bits_in1_7,
  input  [31:0] io_enq_bits_in2_0,
  input  [31:0] io_enq_bits_in2_1,
  input  [31:0] io_enq_bits_in2_2,
  input  [31:0] io_enq_bits_in2_3,
  input  [31:0] io_enq_bits_in2_4,
  input  [31:0] io_enq_bits_in2_5,
  input  [31:0] io_enq_bits_in2_6,
  input  [31:0] io_enq_bits_in2_7,
  input  [31:0] io_enq_bits_in3_0,
  input  [31:0] io_enq_bits_in3_1,
  input  [31:0] io_enq_bits_in3_2,
  input  [31:0] io_enq_bits_in3_3,
  input  [31:0] io_enq_bits_in3_4,
  input  [31:0] io_enq_bits_in3_5,
  input  [31:0] io_enq_bits_in3_6,
  input  [31:0] io_enq_bits_in3_7,
  input         io_enq_bits_mask_0,
  input         io_enq_bits_mask_1,
  input         io_enq_bits_mask_2,
  input         io_enq_bits_mask_3,
  input         io_enq_bits_mask_4,
  input         io_enq_bits_mask_5,
  input         io_enq_bits_mask_6,
  input         io_enq_bits_mask_7,
  input  [31:0] io_enq_bits_ctrl_inst,
  input  [1:0]  io_enq_bits_ctrl_wid,
  input         io_enq_bits_ctrl_fp,
  input  [1:0]  io_enq_bits_ctrl_branch,
  input         io_enq_bits_ctrl_simt_stack,
  input         io_enq_bits_ctrl_simt_stack_op,
  input         io_enq_bits_ctrl_barrier,
  input  [1:0]  io_enq_bits_ctrl_csr,
  input         io_enq_bits_ctrl_reverse,
  input         io_enq_bits_ctrl_isvec,
  input         io_enq_bits_ctrl_mem_unsigned,
  input  [5:0]  io_enq_bits_ctrl_alu_fn,
  input         io_enq_bits_ctrl_mem,
  input  [1:0]  io_enq_bits_ctrl_mem_cmd,
  input  [1:0]  io_enq_bits_ctrl_mop,
  input  [4:0]  io_enq_bits_ctrl_reg_idxw,
  input         io_enq_bits_ctrl_wfd,
  input         io_enq_bits_ctrl_fence,
  input         io_enq_bits_ctrl_sfu,
  input         io_enq_bits_ctrl_readmask,
  input         io_enq_bits_ctrl_writemask,
  input         io_enq_bits_ctrl_wxd,
  input  [31:0] io_enq_bits_ctrl_pc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_in1_0,
  output [31:0] io_deq_bits_in1_1,
  output [31:0] io_deq_bits_in1_2,
  output [31:0] io_deq_bits_in1_3,
  output [31:0] io_deq_bits_in1_4,
  output [31:0] io_deq_bits_in1_5,
  output [31:0] io_deq_bits_in1_6,
  output [31:0] io_deq_bits_in1_7,
  output [31:0] io_deq_bits_in2_0,
  output [31:0] io_deq_bits_in2_1,
  output [31:0] io_deq_bits_in2_2,
  output [31:0] io_deq_bits_in2_3,
  output [31:0] io_deq_bits_in2_4,
  output [31:0] io_deq_bits_in2_5,
  output [31:0] io_deq_bits_in2_6,
  output [31:0] io_deq_bits_in2_7,
  output [31:0] io_deq_bits_in3_0,
  output [31:0] io_deq_bits_in3_1,
  output [31:0] io_deq_bits_in3_2,
  output [31:0] io_deq_bits_in3_3,
  output [31:0] io_deq_bits_in3_4,
  output [31:0] io_deq_bits_in3_5,
  output [31:0] io_deq_bits_in3_6,
  output [31:0] io_deq_bits_in3_7,
  output        io_deq_bits_mask_0,
  output        io_deq_bits_mask_1,
  output        io_deq_bits_mask_2,
  output        io_deq_bits_mask_3,
  output        io_deq_bits_mask_4,
  output        io_deq_bits_mask_5,
  output        io_deq_bits_mask_6,
  output        io_deq_bits_mask_7,
  output [31:0] io_deq_bits_ctrl_inst,
  output [1:0]  io_deq_bits_ctrl_wid,
  output        io_deq_bits_ctrl_fp,
  output [1:0]  io_deq_bits_ctrl_branch,
  output        io_deq_bits_ctrl_simt_stack,
  output        io_deq_bits_ctrl_simt_stack_op,
  output        io_deq_bits_ctrl_barrier,
  output [1:0]  io_deq_bits_ctrl_csr,
  output        io_deq_bits_ctrl_reverse,
  output        io_deq_bits_ctrl_isvec,
  output        io_deq_bits_ctrl_mem_unsigned,
  output [5:0]  io_deq_bits_ctrl_alu_fn,
  output        io_deq_bits_ctrl_mem,
  output [1:0]  io_deq_bits_ctrl_mem_cmd,
  output [1:0]  io_deq_bits_ctrl_mop,
  output [4:0]  io_deq_bits_ctrl_reg_idxw,
  output        io_deq_bits_ctrl_wfd,
  output        io_deq_bits_ctrl_fence,
  output        io_deq_bits_ctrl_sfu,
  output        io_deq_bits_ctrl_readmask,
  output        io_deq_bits_ctrl_writemask,
  output        io_deq_bits_ctrl_wxd,
  output [31:0] io_deq_bits_ctrl_pc
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_55;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_in1_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in3_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in3_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in3_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in3_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in3_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in3_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in3_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_ctrl_inst [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_inst_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_inst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_ctrl_inst_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_ctrl_inst_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_inst_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_inst_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_inst_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_ctrl_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_fp [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_ctrl_branch [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_branch_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_branch_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_branch_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_branch_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_branch_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_branch_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_branch_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_simt_stack [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_simt_stack_op [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_simt_stack_op_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_barrier [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_barrier_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_ctrl_csr [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_csr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_csr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_csr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_csr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_csr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_csr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_csr_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_reverse [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_isvec [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_mem_unsigned [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_unsigned_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] ram_ctrl_alu_fn [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [5:0] ram_ctrl_alu_fn_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_ctrl_alu_fn_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_mem [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_ctrl_mem_cmd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_cmd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_cmd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_mem_cmd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_mem_cmd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_cmd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_cmd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mem_cmd_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_ctrl_mop [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mop_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mop_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_mop_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_mop_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mop_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mop_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_mop_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_ctrl_reg_idxw [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wfd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_fence [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fence_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_sfu [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_sfu_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_readmask [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_readmask_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_writemask [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_writemask_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wxd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_ctrl_pc [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_pc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_pc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_ctrl_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_ctrl_pc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_pc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_pc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_pc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_in1_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_0_io_deq_bits_MPORT_data = ram_in1_0[ram_in1_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_0_MPORT_data = io_enq_bits_in1_0;
  assign ram_in1_0_MPORT_addr = 1'h0;
  assign ram_in1_0_MPORT_mask = 1'h1;
  assign ram_in1_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_1_io_deq_bits_MPORT_data = ram_in1_1[ram_in1_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_1_MPORT_data = io_enq_bits_in1_1;
  assign ram_in1_1_MPORT_addr = 1'h0;
  assign ram_in1_1_MPORT_mask = 1'h1;
  assign ram_in1_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_2_io_deq_bits_MPORT_data = ram_in1_2[ram_in1_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_2_MPORT_data = io_enq_bits_in1_2;
  assign ram_in1_2_MPORT_addr = 1'h0;
  assign ram_in1_2_MPORT_mask = 1'h1;
  assign ram_in1_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_3_io_deq_bits_MPORT_data = ram_in1_3[ram_in1_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_3_MPORT_data = io_enq_bits_in1_3;
  assign ram_in1_3_MPORT_addr = 1'h0;
  assign ram_in1_3_MPORT_mask = 1'h1;
  assign ram_in1_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_4_io_deq_bits_MPORT_data = ram_in1_4[ram_in1_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_4_MPORT_data = io_enq_bits_in1_4;
  assign ram_in1_4_MPORT_addr = 1'h0;
  assign ram_in1_4_MPORT_mask = 1'h1;
  assign ram_in1_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_5_io_deq_bits_MPORT_data = ram_in1_5[ram_in1_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_5_MPORT_data = io_enq_bits_in1_5;
  assign ram_in1_5_MPORT_addr = 1'h0;
  assign ram_in1_5_MPORT_mask = 1'h1;
  assign ram_in1_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_6_io_deq_bits_MPORT_data = ram_in1_6[ram_in1_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_6_MPORT_data = io_enq_bits_in1_6;
  assign ram_in1_6_MPORT_addr = 1'h0;
  assign ram_in1_6_MPORT_mask = 1'h1;
  assign ram_in1_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_7_io_deq_bits_MPORT_data = ram_in1_7[ram_in1_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_7_MPORT_data = io_enq_bits_in1_7;
  assign ram_in1_7_MPORT_addr = 1'h0;
  assign ram_in1_7_MPORT_mask = 1'h1;
  assign ram_in1_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_0_io_deq_bits_MPORT_data = ram_in2_0[ram_in2_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_0_MPORT_data = io_enq_bits_in2_0;
  assign ram_in2_0_MPORT_addr = 1'h0;
  assign ram_in2_0_MPORT_mask = 1'h1;
  assign ram_in2_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_1_io_deq_bits_MPORT_data = ram_in2_1[ram_in2_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_1_MPORT_data = io_enq_bits_in2_1;
  assign ram_in2_1_MPORT_addr = 1'h0;
  assign ram_in2_1_MPORT_mask = 1'h1;
  assign ram_in2_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_2_io_deq_bits_MPORT_data = ram_in2_2[ram_in2_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_2_MPORT_data = io_enq_bits_in2_2;
  assign ram_in2_2_MPORT_addr = 1'h0;
  assign ram_in2_2_MPORT_mask = 1'h1;
  assign ram_in2_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_3_io_deq_bits_MPORT_data = ram_in2_3[ram_in2_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_3_MPORT_data = io_enq_bits_in2_3;
  assign ram_in2_3_MPORT_addr = 1'h0;
  assign ram_in2_3_MPORT_mask = 1'h1;
  assign ram_in2_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_4_io_deq_bits_MPORT_data = ram_in2_4[ram_in2_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_4_MPORT_data = io_enq_bits_in2_4;
  assign ram_in2_4_MPORT_addr = 1'h0;
  assign ram_in2_4_MPORT_mask = 1'h1;
  assign ram_in2_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_5_io_deq_bits_MPORT_data = ram_in2_5[ram_in2_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_5_MPORT_data = io_enq_bits_in2_5;
  assign ram_in2_5_MPORT_addr = 1'h0;
  assign ram_in2_5_MPORT_mask = 1'h1;
  assign ram_in2_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_6_io_deq_bits_MPORT_data = ram_in2_6[ram_in2_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_6_MPORT_data = io_enq_bits_in2_6;
  assign ram_in2_6_MPORT_addr = 1'h0;
  assign ram_in2_6_MPORT_mask = 1'h1;
  assign ram_in2_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_7_io_deq_bits_MPORT_data = ram_in2_7[ram_in2_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_7_MPORT_data = io_enq_bits_in2_7;
  assign ram_in2_7_MPORT_addr = 1'h0;
  assign ram_in2_7_MPORT_mask = 1'h1;
  assign ram_in2_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_0_io_deq_bits_MPORT_data = ram_in3_0[ram_in3_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_0_MPORT_data = io_enq_bits_in3_0;
  assign ram_in3_0_MPORT_addr = 1'h0;
  assign ram_in3_0_MPORT_mask = 1'h1;
  assign ram_in3_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_1_io_deq_bits_MPORT_data = ram_in3_1[ram_in3_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_1_MPORT_data = io_enq_bits_in3_1;
  assign ram_in3_1_MPORT_addr = 1'h0;
  assign ram_in3_1_MPORT_mask = 1'h1;
  assign ram_in3_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_2_io_deq_bits_MPORT_data = ram_in3_2[ram_in3_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_2_MPORT_data = io_enq_bits_in3_2;
  assign ram_in3_2_MPORT_addr = 1'h0;
  assign ram_in3_2_MPORT_mask = 1'h1;
  assign ram_in3_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_3_io_deq_bits_MPORT_data = ram_in3_3[ram_in3_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_3_MPORT_data = io_enq_bits_in3_3;
  assign ram_in3_3_MPORT_addr = 1'h0;
  assign ram_in3_3_MPORT_mask = 1'h1;
  assign ram_in3_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_4_io_deq_bits_MPORT_data = ram_in3_4[ram_in3_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_4_MPORT_data = io_enq_bits_in3_4;
  assign ram_in3_4_MPORT_addr = 1'h0;
  assign ram_in3_4_MPORT_mask = 1'h1;
  assign ram_in3_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_5_io_deq_bits_MPORT_data = ram_in3_5[ram_in3_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_5_MPORT_data = io_enq_bits_in3_5;
  assign ram_in3_5_MPORT_addr = 1'h0;
  assign ram_in3_5_MPORT_mask = 1'h1;
  assign ram_in3_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_6_io_deq_bits_MPORT_data = ram_in3_6[ram_in3_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_6_MPORT_data = io_enq_bits_in3_6;
  assign ram_in3_6_MPORT_addr = 1'h0;
  assign ram_in3_6_MPORT_mask = 1'h1;
  assign ram_in3_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in3_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in3_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in3_7_io_deq_bits_MPORT_data = ram_in3_7[ram_in3_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in3_7_MPORT_data = io_enq_bits_in3_7;
  assign ram_in3_7_MPORT_addr = 1'h0;
  assign ram_in3_7_MPORT_mask = 1'h1;
  assign ram_in3_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_0_io_deq_bits_MPORT_data = ram_mask_0[ram_mask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_0_MPORT_data = io_enq_bits_mask_0;
  assign ram_mask_0_MPORT_addr = 1'h0;
  assign ram_mask_0_MPORT_mask = 1'h1;
  assign ram_mask_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_1_io_deq_bits_MPORT_data = ram_mask_1[ram_mask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_1_MPORT_data = io_enq_bits_mask_1;
  assign ram_mask_1_MPORT_addr = 1'h0;
  assign ram_mask_1_MPORT_mask = 1'h1;
  assign ram_mask_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_2_io_deq_bits_MPORT_data = ram_mask_2[ram_mask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_2_MPORT_data = io_enq_bits_mask_2;
  assign ram_mask_2_MPORT_addr = 1'h0;
  assign ram_mask_2_MPORT_mask = 1'h1;
  assign ram_mask_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_3_io_deq_bits_MPORT_data = ram_mask_3[ram_mask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_3_MPORT_data = io_enq_bits_mask_3;
  assign ram_mask_3_MPORT_addr = 1'h0;
  assign ram_mask_3_MPORT_mask = 1'h1;
  assign ram_mask_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_4_io_deq_bits_MPORT_data = ram_mask_4[ram_mask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_4_MPORT_data = io_enq_bits_mask_4;
  assign ram_mask_4_MPORT_addr = 1'h0;
  assign ram_mask_4_MPORT_mask = 1'h1;
  assign ram_mask_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_5_io_deq_bits_MPORT_data = ram_mask_5[ram_mask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_5_MPORT_data = io_enq_bits_mask_5;
  assign ram_mask_5_MPORT_addr = 1'h0;
  assign ram_mask_5_MPORT_mask = 1'h1;
  assign ram_mask_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_6_io_deq_bits_MPORT_data = ram_mask_6[ram_mask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_6_MPORT_data = io_enq_bits_mask_6;
  assign ram_mask_6_MPORT_addr = 1'h0;
  assign ram_mask_6_MPORT_mask = 1'h1;
  assign ram_mask_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_7_io_deq_bits_MPORT_data = ram_mask_7[ram_mask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_7_MPORT_data = io_enq_bits_mask_7;
  assign ram_mask_7_MPORT_addr = 1'h0;
  assign ram_mask_7_MPORT_mask = 1'h1;
  assign ram_mask_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_inst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_inst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_inst_io_deq_bits_MPORT_data = ram_ctrl_inst[ram_ctrl_inst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_inst_MPORT_data = io_enq_bits_ctrl_inst;
  assign ram_ctrl_inst_MPORT_addr = 1'h0;
  assign ram_ctrl_inst_MPORT_mask = 1'h1;
  assign ram_ctrl_inst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wid_io_deq_bits_MPORT_data = ram_ctrl_wid[ram_ctrl_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wid_MPORT_data = io_enq_bits_ctrl_wid;
  assign ram_ctrl_wid_MPORT_addr = 1'h0;
  assign ram_ctrl_wid_MPORT_mask = 1'h1;
  assign ram_ctrl_wid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_fp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_fp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_fp_io_deq_bits_MPORT_data = ram_ctrl_fp[ram_ctrl_fp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_fp_MPORT_data = io_enq_bits_ctrl_fp;
  assign ram_ctrl_fp_MPORT_addr = 1'h0;
  assign ram_ctrl_fp_MPORT_mask = 1'h1;
  assign ram_ctrl_fp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_branch_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_branch_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_branch_io_deq_bits_MPORT_data = ram_ctrl_branch[ram_ctrl_branch_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_branch_MPORT_data = io_enq_bits_ctrl_branch;
  assign ram_ctrl_branch_MPORT_addr = 1'h0;
  assign ram_ctrl_branch_MPORT_mask = 1'h1;
  assign ram_ctrl_branch_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_simt_stack_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_simt_stack_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_simt_stack_io_deq_bits_MPORT_data = ram_ctrl_simt_stack[ram_ctrl_simt_stack_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_simt_stack_MPORT_data = io_enq_bits_ctrl_simt_stack;
  assign ram_ctrl_simt_stack_MPORT_addr = 1'h0;
  assign ram_ctrl_simt_stack_MPORT_mask = 1'h1;
  assign ram_ctrl_simt_stack_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_simt_stack_op_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_simt_stack_op_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_simt_stack_op_io_deq_bits_MPORT_data =
    ram_ctrl_simt_stack_op[ram_ctrl_simt_stack_op_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_simt_stack_op_MPORT_data = io_enq_bits_ctrl_simt_stack_op;
  assign ram_ctrl_simt_stack_op_MPORT_addr = 1'h0;
  assign ram_ctrl_simt_stack_op_MPORT_mask = 1'h1;
  assign ram_ctrl_simt_stack_op_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_barrier_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_barrier_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_barrier_io_deq_bits_MPORT_data = ram_ctrl_barrier[ram_ctrl_barrier_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_barrier_MPORT_data = io_enq_bits_ctrl_barrier;
  assign ram_ctrl_barrier_MPORT_addr = 1'h0;
  assign ram_ctrl_barrier_MPORT_mask = 1'h1;
  assign ram_ctrl_barrier_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_csr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_csr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_csr_io_deq_bits_MPORT_data = ram_ctrl_csr[ram_ctrl_csr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_csr_MPORT_data = io_enq_bits_ctrl_csr;
  assign ram_ctrl_csr_MPORT_addr = 1'h0;
  assign ram_ctrl_csr_MPORT_mask = 1'h1;
  assign ram_ctrl_csr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_reverse_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_reverse_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_reverse_io_deq_bits_MPORT_data = ram_ctrl_reverse[ram_ctrl_reverse_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_reverse_MPORT_data = io_enq_bits_ctrl_reverse;
  assign ram_ctrl_reverse_MPORT_addr = 1'h0;
  assign ram_ctrl_reverse_MPORT_mask = 1'h1;
  assign ram_ctrl_reverse_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_isvec_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_isvec_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_isvec_io_deq_bits_MPORT_data = ram_ctrl_isvec[ram_ctrl_isvec_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_isvec_MPORT_data = io_enq_bits_ctrl_isvec;
  assign ram_ctrl_isvec_MPORT_addr = 1'h0;
  assign ram_ctrl_isvec_MPORT_mask = 1'h1;
  assign ram_ctrl_isvec_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_mem_unsigned_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_mem_unsigned_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_mem_unsigned_io_deq_bits_MPORT_data =
    ram_ctrl_mem_unsigned[ram_ctrl_mem_unsigned_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_mem_unsigned_MPORT_data = io_enq_bits_ctrl_mem_unsigned;
  assign ram_ctrl_mem_unsigned_MPORT_addr = 1'h0;
  assign ram_ctrl_mem_unsigned_MPORT_mask = 1'h1;
  assign ram_ctrl_mem_unsigned_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_alu_fn_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_alu_fn_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_alu_fn_io_deq_bits_MPORT_data = ram_ctrl_alu_fn[ram_ctrl_alu_fn_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_alu_fn_MPORT_data = io_enq_bits_ctrl_alu_fn;
  assign ram_ctrl_alu_fn_MPORT_addr = 1'h0;
  assign ram_ctrl_alu_fn_MPORT_mask = 1'h1;
  assign ram_ctrl_alu_fn_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_mem_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_mem_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_mem_io_deq_bits_MPORT_data = ram_ctrl_mem[ram_ctrl_mem_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_mem_MPORT_data = io_enq_bits_ctrl_mem;
  assign ram_ctrl_mem_MPORT_addr = 1'h0;
  assign ram_ctrl_mem_MPORT_mask = 1'h1;
  assign ram_ctrl_mem_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_mem_cmd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_mem_cmd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_mem_cmd_io_deq_bits_MPORT_data = ram_ctrl_mem_cmd[ram_ctrl_mem_cmd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_mem_cmd_MPORT_data = io_enq_bits_ctrl_mem_cmd;
  assign ram_ctrl_mem_cmd_MPORT_addr = 1'h0;
  assign ram_ctrl_mem_cmd_MPORT_mask = 1'h1;
  assign ram_ctrl_mem_cmd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_mop_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_mop_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_mop_io_deq_bits_MPORT_data = ram_ctrl_mop[ram_ctrl_mop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_mop_MPORT_data = io_enq_bits_ctrl_mop;
  assign ram_ctrl_mop_MPORT_addr = 1'h0;
  assign ram_ctrl_mop_MPORT_mask = 1'h1;
  assign ram_ctrl_mop_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_data = ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_reg_idxw_MPORT_data = io_enq_bits_ctrl_reg_idxw;
  assign ram_ctrl_reg_idxw_MPORT_addr = 1'h0;
  assign ram_ctrl_reg_idxw_MPORT_mask = 1'h1;
  assign ram_ctrl_reg_idxw_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_data = ram_ctrl_wfd[ram_ctrl_wfd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wfd_MPORT_data = io_enq_bits_ctrl_wfd;
  assign ram_ctrl_wfd_MPORT_addr = 1'h0;
  assign ram_ctrl_wfd_MPORT_mask = 1'h1;
  assign ram_ctrl_wfd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_fence_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_fence_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_fence_io_deq_bits_MPORT_data = ram_ctrl_fence[ram_ctrl_fence_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_fence_MPORT_data = io_enq_bits_ctrl_fence;
  assign ram_ctrl_fence_MPORT_addr = 1'h0;
  assign ram_ctrl_fence_MPORT_mask = 1'h1;
  assign ram_ctrl_fence_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_sfu_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_sfu_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_sfu_io_deq_bits_MPORT_data = ram_ctrl_sfu[ram_ctrl_sfu_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_sfu_MPORT_data = io_enq_bits_ctrl_sfu;
  assign ram_ctrl_sfu_MPORT_addr = 1'h0;
  assign ram_ctrl_sfu_MPORT_mask = 1'h1;
  assign ram_ctrl_sfu_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_readmask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_readmask_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_readmask_io_deq_bits_MPORT_data = ram_ctrl_readmask[ram_ctrl_readmask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_readmask_MPORT_data = io_enq_bits_ctrl_readmask;
  assign ram_ctrl_readmask_MPORT_addr = 1'h0;
  assign ram_ctrl_readmask_MPORT_mask = 1'h1;
  assign ram_ctrl_readmask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_writemask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_writemask_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_writemask_io_deq_bits_MPORT_data = ram_ctrl_writemask[ram_ctrl_writemask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_writemask_MPORT_data = io_enq_bits_ctrl_writemask;
  assign ram_ctrl_writemask_MPORT_addr = 1'h0;
  assign ram_ctrl_writemask_MPORT_mask = 1'h1;
  assign ram_ctrl_writemask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_data = ram_ctrl_wxd[ram_ctrl_wxd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wxd_MPORT_data = io_enq_bits_ctrl_wxd;
  assign ram_ctrl_wxd_MPORT_addr = 1'h0;
  assign ram_ctrl_wxd_MPORT_mask = 1'h1;
  assign ram_ctrl_wxd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_pc_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_pc_io_deq_bits_MPORT_data = ram_ctrl_pc[ram_ctrl_pc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_pc_MPORT_data = io_enq_bits_ctrl_pc;
  assign ram_ctrl_pc_MPORT_addr = 1'h0;
  assign ram_ctrl_pc_MPORT_mask = 1'h1;
  assign ram_ctrl_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_in1_0 = ram_in1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_1 = ram_in1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_2 = ram_in1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_3 = ram_in1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_4 = ram_in1_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_5 = ram_in1_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_6 = ram_in1_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_7 = ram_in1_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_0 = ram_in2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_1 = ram_in2_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_2 = ram_in2_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_3 = ram_in2_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_4 = ram_in2_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_5 = ram_in2_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_6 = ram_in2_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_7 = ram_in2_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_0 = ram_in3_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_1 = ram_in3_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_2 = ram_in3_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_3 = ram_in3_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_4 = ram_in3_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_5 = ram_in3_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_6 = ram_in3_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in3_7 = ram_in3_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_0 = ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_1 = ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_2 = ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_3 = ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_4 = ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_5 = ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_6 = ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_7 = ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_inst = ram_ctrl_inst_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_wid = ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_fp = ram_ctrl_fp_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_branch = ram_ctrl_branch_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_simt_stack = ram_ctrl_simt_stack_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_simt_stack_op = ram_ctrl_simt_stack_op_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_barrier = ram_ctrl_barrier_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_csr = ram_ctrl_csr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_reverse = ram_ctrl_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_isvec = ram_ctrl_isvec_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_mem_unsigned = ram_ctrl_mem_unsigned_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_alu_fn = ram_ctrl_alu_fn_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_mem = ram_ctrl_mem_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_mem_cmd = ram_ctrl_mem_cmd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_mop = ram_ctrl_mop_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_reg_idxw = ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_wfd = ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_fence = ram_ctrl_fence_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_sfu = ram_ctrl_sfu_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_readmask = ram_ctrl_readmask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_writemask = ram_ctrl_writemask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_wxd = ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_pc = ram_ctrl_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_in1_0_MPORT_en & ram_in1_0_MPORT_mask) begin
      ram_in1_0[ram_in1_0_MPORT_addr] <= ram_in1_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_1_MPORT_en & ram_in1_1_MPORT_mask) begin
      ram_in1_1[ram_in1_1_MPORT_addr] <= ram_in1_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_2_MPORT_en & ram_in1_2_MPORT_mask) begin
      ram_in1_2[ram_in1_2_MPORT_addr] <= ram_in1_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_3_MPORT_en & ram_in1_3_MPORT_mask) begin
      ram_in1_3[ram_in1_3_MPORT_addr] <= ram_in1_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_4_MPORT_en & ram_in1_4_MPORT_mask) begin
      ram_in1_4[ram_in1_4_MPORT_addr] <= ram_in1_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_5_MPORT_en & ram_in1_5_MPORT_mask) begin
      ram_in1_5[ram_in1_5_MPORT_addr] <= ram_in1_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_6_MPORT_en & ram_in1_6_MPORT_mask) begin
      ram_in1_6[ram_in1_6_MPORT_addr] <= ram_in1_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_7_MPORT_en & ram_in1_7_MPORT_mask) begin
      ram_in1_7[ram_in1_7_MPORT_addr] <= ram_in1_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_0_MPORT_en & ram_in2_0_MPORT_mask) begin
      ram_in2_0[ram_in2_0_MPORT_addr] <= ram_in2_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_1_MPORT_en & ram_in2_1_MPORT_mask) begin
      ram_in2_1[ram_in2_1_MPORT_addr] <= ram_in2_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_2_MPORT_en & ram_in2_2_MPORT_mask) begin
      ram_in2_2[ram_in2_2_MPORT_addr] <= ram_in2_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_3_MPORT_en & ram_in2_3_MPORT_mask) begin
      ram_in2_3[ram_in2_3_MPORT_addr] <= ram_in2_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_4_MPORT_en & ram_in2_4_MPORT_mask) begin
      ram_in2_4[ram_in2_4_MPORT_addr] <= ram_in2_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_5_MPORT_en & ram_in2_5_MPORT_mask) begin
      ram_in2_5[ram_in2_5_MPORT_addr] <= ram_in2_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_6_MPORT_en & ram_in2_6_MPORT_mask) begin
      ram_in2_6[ram_in2_6_MPORT_addr] <= ram_in2_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_7_MPORT_en & ram_in2_7_MPORT_mask) begin
      ram_in2_7[ram_in2_7_MPORT_addr] <= ram_in2_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_0_MPORT_en & ram_in3_0_MPORT_mask) begin
      ram_in3_0[ram_in3_0_MPORT_addr] <= ram_in3_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_1_MPORT_en & ram_in3_1_MPORT_mask) begin
      ram_in3_1[ram_in3_1_MPORT_addr] <= ram_in3_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_2_MPORT_en & ram_in3_2_MPORT_mask) begin
      ram_in3_2[ram_in3_2_MPORT_addr] <= ram_in3_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_3_MPORT_en & ram_in3_3_MPORT_mask) begin
      ram_in3_3[ram_in3_3_MPORT_addr] <= ram_in3_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_4_MPORT_en & ram_in3_4_MPORT_mask) begin
      ram_in3_4[ram_in3_4_MPORT_addr] <= ram_in3_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_5_MPORT_en & ram_in3_5_MPORT_mask) begin
      ram_in3_5[ram_in3_5_MPORT_addr] <= ram_in3_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_6_MPORT_en & ram_in3_6_MPORT_mask) begin
      ram_in3_6[ram_in3_6_MPORT_addr] <= ram_in3_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in3_7_MPORT_en & ram_in3_7_MPORT_mask) begin
      ram_in3_7[ram_in3_7_MPORT_addr] <= ram_in3_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_0_MPORT_en & ram_mask_0_MPORT_mask) begin
      ram_mask_0[ram_mask_0_MPORT_addr] <= ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_1_MPORT_en & ram_mask_1_MPORT_mask) begin
      ram_mask_1[ram_mask_1_MPORT_addr] <= ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_2_MPORT_en & ram_mask_2_MPORT_mask) begin
      ram_mask_2[ram_mask_2_MPORT_addr] <= ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_3_MPORT_en & ram_mask_3_MPORT_mask) begin
      ram_mask_3[ram_mask_3_MPORT_addr] <= ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_4_MPORT_en & ram_mask_4_MPORT_mask) begin
      ram_mask_4[ram_mask_4_MPORT_addr] <= ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_5_MPORT_en & ram_mask_5_MPORT_mask) begin
      ram_mask_5[ram_mask_5_MPORT_addr] <= ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_6_MPORT_en & ram_mask_6_MPORT_mask) begin
      ram_mask_6[ram_mask_6_MPORT_addr] <= ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_7_MPORT_en & ram_mask_7_MPORT_mask) begin
      ram_mask_7[ram_mask_7_MPORT_addr] <= ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_inst_MPORT_en & ram_ctrl_inst_MPORT_mask) begin
      ram_ctrl_inst[ram_ctrl_inst_MPORT_addr] <= ram_ctrl_inst_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wid_MPORT_en & ram_ctrl_wid_MPORT_mask) begin
      ram_ctrl_wid[ram_ctrl_wid_MPORT_addr] <= ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_fp_MPORT_en & ram_ctrl_fp_MPORT_mask) begin
      ram_ctrl_fp[ram_ctrl_fp_MPORT_addr] <= ram_ctrl_fp_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_branch_MPORT_en & ram_ctrl_branch_MPORT_mask) begin
      ram_ctrl_branch[ram_ctrl_branch_MPORT_addr] <= ram_ctrl_branch_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_simt_stack_MPORT_en & ram_ctrl_simt_stack_MPORT_mask) begin
      ram_ctrl_simt_stack[ram_ctrl_simt_stack_MPORT_addr] <= ram_ctrl_simt_stack_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_simt_stack_op_MPORT_en & ram_ctrl_simt_stack_op_MPORT_mask) begin
      ram_ctrl_simt_stack_op[ram_ctrl_simt_stack_op_MPORT_addr] <= ram_ctrl_simt_stack_op_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_barrier_MPORT_en & ram_ctrl_barrier_MPORT_mask) begin
      ram_ctrl_barrier[ram_ctrl_barrier_MPORT_addr] <= ram_ctrl_barrier_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_csr_MPORT_en & ram_ctrl_csr_MPORT_mask) begin
      ram_ctrl_csr[ram_ctrl_csr_MPORT_addr] <= ram_ctrl_csr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_reverse_MPORT_en & ram_ctrl_reverse_MPORT_mask) begin
      ram_ctrl_reverse[ram_ctrl_reverse_MPORT_addr] <= ram_ctrl_reverse_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_isvec_MPORT_en & ram_ctrl_isvec_MPORT_mask) begin
      ram_ctrl_isvec[ram_ctrl_isvec_MPORT_addr] <= ram_ctrl_isvec_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_mem_unsigned_MPORT_en & ram_ctrl_mem_unsigned_MPORT_mask) begin
      ram_ctrl_mem_unsigned[ram_ctrl_mem_unsigned_MPORT_addr] <= ram_ctrl_mem_unsigned_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_alu_fn_MPORT_en & ram_ctrl_alu_fn_MPORT_mask) begin
      ram_ctrl_alu_fn[ram_ctrl_alu_fn_MPORT_addr] <= ram_ctrl_alu_fn_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_mem_MPORT_en & ram_ctrl_mem_MPORT_mask) begin
      ram_ctrl_mem[ram_ctrl_mem_MPORT_addr] <= ram_ctrl_mem_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_mem_cmd_MPORT_en & ram_ctrl_mem_cmd_MPORT_mask) begin
      ram_ctrl_mem_cmd[ram_ctrl_mem_cmd_MPORT_addr] <= ram_ctrl_mem_cmd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_mop_MPORT_en & ram_ctrl_mop_MPORT_mask) begin
      ram_ctrl_mop[ram_ctrl_mop_MPORT_addr] <= ram_ctrl_mop_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_reg_idxw_MPORT_en & ram_ctrl_reg_idxw_MPORT_mask) begin
      ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_MPORT_addr] <= ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wfd_MPORT_en & ram_ctrl_wfd_MPORT_mask) begin
      ram_ctrl_wfd[ram_ctrl_wfd_MPORT_addr] <= ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_fence_MPORT_en & ram_ctrl_fence_MPORT_mask) begin
      ram_ctrl_fence[ram_ctrl_fence_MPORT_addr] <= ram_ctrl_fence_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_sfu_MPORT_en & ram_ctrl_sfu_MPORT_mask) begin
      ram_ctrl_sfu[ram_ctrl_sfu_MPORT_addr] <= ram_ctrl_sfu_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_readmask_MPORT_en & ram_ctrl_readmask_MPORT_mask) begin
      ram_ctrl_readmask[ram_ctrl_readmask_MPORT_addr] <= ram_ctrl_readmask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_writemask_MPORT_en & ram_ctrl_writemask_MPORT_mask) begin
      ram_ctrl_writemask[ram_ctrl_writemask_MPORT_addr] <= ram_ctrl_writemask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wxd_MPORT_en & ram_ctrl_wxd_MPORT_mask) begin
      ram_ctrl_wxd[ram_ctrl_wxd_MPORT_addr] <= ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_pc_MPORT_en & ram_ctrl_pc_MPORT_mask) begin
      ram_ctrl_pc[ram_ctrl_pc_MPORT_addr] <= ram_ctrl_pc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_0[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_1[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_2[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_3[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_4[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_5[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_6[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_7[initvar] = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_0[initvar] = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_1[initvar] = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_2[initvar] = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_3[initvar] = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_4[initvar] = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_5[initvar] = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_6[initvar] = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_7[initvar] = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_0[initvar] = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_1[initvar] = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_2[initvar] = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_3[initvar] = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_4[initvar] = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_5[initvar] = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_6[initvar] = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in3_7[initvar] = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_0[initvar] = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_1[initvar] = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_2[initvar] = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_3[initvar] = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_4[initvar] = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_5[initvar] = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_6[initvar] = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_7[initvar] = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_inst[initvar] = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wid[initvar] = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_fp[initvar] = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_branch[initvar] = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_simt_stack[initvar] = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_simt_stack_op[initvar] = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_barrier[initvar] = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_csr[initvar] = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_reverse[initvar] = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_isvec[initvar] = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_mem_unsigned[initvar] = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_alu_fn[initvar] = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_mem[initvar] = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_mem_cmd[initvar] = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_mop[initvar] = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_reg_idxw[initvar] = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wfd[initvar] = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_fence[initvar] = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_sfu[initvar] = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_readmask[initvar] = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_writemask[initvar] = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wxd[initvar] = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_pc[initvar] = _RAND_54[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  maybe_full = _RAND_55[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AddrCalculate(
  input         clock,
  input         reset,
  output        io_from_fifo_ready,
  input         io_from_fifo_valid,
  input  [31:0] io_from_fifo_bits_in1_0,
  input  [31:0] io_from_fifo_bits_in1_1,
  input  [31:0] io_from_fifo_bits_in1_2,
  input  [31:0] io_from_fifo_bits_in1_3,
  input  [31:0] io_from_fifo_bits_in1_4,
  input  [31:0] io_from_fifo_bits_in1_5,
  input  [31:0] io_from_fifo_bits_in1_6,
  input  [31:0] io_from_fifo_bits_in1_7,
  input  [31:0] io_from_fifo_bits_in2_0,
  input  [31:0] io_from_fifo_bits_in2_1,
  input  [31:0] io_from_fifo_bits_in2_2,
  input  [31:0] io_from_fifo_bits_in2_3,
  input  [31:0] io_from_fifo_bits_in2_4,
  input  [31:0] io_from_fifo_bits_in2_5,
  input  [31:0] io_from_fifo_bits_in2_6,
  input  [31:0] io_from_fifo_bits_in2_7,
  input  [31:0] io_from_fifo_bits_in3_0,
  input  [31:0] io_from_fifo_bits_in3_1,
  input  [31:0] io_from_fifo_bits_in3_2,
  input  [31:0] io_from_fifo_bits_in3_3,
  input  [31:0] io_from_fifo_bits_in3_4,
  input  [31:0] io_from_fifo_bits_in3_5,
  input  [31:0] io_from_fifo_bits_in3_6,
  input  [31:0] io_from_fifo_bits_in3_7,
  input         io_from_fifo_bits_mask_0,
  input         io_from_fifo_bits_mask_1,
  input         io_from_fifo_bits_mask_2,
  input         io_from_fifo_bits_mask_3,
  input         io_from_fifo_bits_mask_4,
  input         io_from_fifo_bits_mask_5,
  input         io_from_fifo_bits_mask_6,
  input         io_from_fifo_bits_mask_7,
  input  [1:0]  io_from_fifo_bits_ctrl_wid,
  input         io_from_fifo_bits_ctrl_isvec,
  input         io_from_fifo_bits_ctrl_mem_unsigned,
  input  [1:0]  io_from_fifo_bits_ctrl_mem_cmd,
  input  [1:0]  io_from_fifo_bits_ctrl_mop,
  input  [4:0]  io_from_fifo_bits_ctrl_reg_idxw,
  input         io_from_fifo_bits_ctrl_wfd,
  input         io_from_fifo_bits_ctrl_wxd,
  input         io_to_mshr_ready,
  output        io_to_mshr_valid,
  output [1:0]  io_to_mshr_bits_tag_warp_id,
  output        io_to_mshr_bits_tag_wfd,
  output        io_to_mshr_bits_tag_wxd,
  output [4:0]  io_to_mshr_bits_tag_reg_idxw,
  output        io_to_mshr_bits_tag_mask_0,
  output        io_to_mshr_bits_tag_mask_1,
  output        io_to_mshr_bits_tag_mask_2,
  output        io_to_mshr_bits_tag_mask_3,
  output        io_to_mshr_bits_tag_mask_4,
  output        io_to_mshr_bits_tag_mask_5,
  output        io_to_mshr_bits_tag_mask_6,
  output        io_to_mshr_bits_tag_mask_7,
  output        io_to_mshr_bits_tag_unsigned,
  output        io_to_mshr_bits_tag_isvec,
  output        io_to_mshr_bits_tag_isWrite,
  input  [1:0]  io_idx_entry,
  input         io_to_dcache_ready,
  output        io_to_dcache_valid,
  output [1:0]  io_to_dcache_bits_instrId,
  output        io_to_dcache_bits_isWrite,
  output [21:0] io_to_dcache_bits_tag,
  output [4:0]  io_to_dcache_bits_setIdx,
  output        io_to_dcache_bits_perLaneAddr_0_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_0_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_1_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_1_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_2_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_2_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_3_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_3_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_4_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_4_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_5_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_5_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_6_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_6_blockOffset,
  output        io_to_dcache_bits_perLaneAddr_7_activeMask,
  output [2:0]  io_to_dcache_bits_perLaneAddr_7_blockOffset,
  output [31:0] io_to_dcache_bits_data_0,
  output [31:0] io_to_dcache_bits_data_1,
  output [31:0] io_to_dcache_bits_data_2,
  output [31:0] io_to_dcache_bits_data_3,
  output [31:0] io_to_dcache_bits_data_4,
  output [31:0] io_to_dcache_bits_data_5,
  output [31:0] io_to_dcache_bits_data_6,
  output [31:0] io_to_dcache_bits_data_7,
  input         io_to_shared_ready,
  output        io_to_shared_valid,
  output [1:0]  io_to_shared_bits_instrId,
  output        io_to_shared_bits_isWrite,
  output [4:0]  io_to_shared_bits_setIdx,
  output        io_to_shared_bits_perLaneAddr_0_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_0_blockOffset,
  output        io_to_shared_bits_perLaneAddr_1_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_1_blockOffset,
  output        io_to_shared_bits_perLaneAddr_2_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_2_blockOffset,
  output        io_to_shared_bits_perLaneAddr_3_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_3_blockOffset,
  output        io_to_shared_bits_perLaneAddr_4_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_4_blockOffset,
  output        io_to_shared_bits_perLaneAddr_5_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_5_blockOffset,
  output        io_to_shared_bits_perLaneAddr_6_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_6_blockOffset,
  output        io_to_shared_bits_perLaneAddr_7_activeMask,
  output [2:0]  io_to_shared_bits_perLaneAddr_7_blockOffset,
  output [31:0] io_to_shared_bits_data_0,
  output [31:0] io_to_shared_bits_data_1,
  output [31:0] io_to_shared_bits_data_2,
  output [31:0] io_to_shared_bits_data_3,
  output [31:0] io_to_shared_bits_data_4,
  output [31:0] io_to_shared_bits_data_5,
  output [31:0] io_to_shared_bits_data_6,
  output [31:0] io_to_shared_bits_data_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[LSU.scala 131:22]
  reg [31:0] reg_save_in1_0; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_1; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_2; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_3; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_4; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_5; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_6; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in1_7; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_0; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_1; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_2; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_3; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_4; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_5; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_6; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in2_7; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_0; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_1; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_2; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_3; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_4; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_5; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_6; // @[LSU.scala 133:21]
  reg [31:0] reg_save_in3_7; // @[LSU.scala 133:21]
  reg  reg_save_mask_0; // @[LSU.scala 133:21]
  reg  reg_save_mask_1; // @[LSU.scala 133:21]
  reg  reg_save_mask_2; // @[LSU.scala 133:21]
  reg  reg_save_mask_3; // @[LSU.scala 133:21]
  reg  reg_save_mask_4; // @[LSU.scala 133:21]
  reg  reg_save_mask_5; // @[LSU.scala 133:21]
  reg  reg_save_mask_6; // @[LSU.scala 133:21]
  reg  reg_save_mask_7; // @[LSU.scala 133:21]
  reg [1:0] reg_save_ctrl_wid; // @[LSU.scala 133:21]
  reg  reg_save_ctrl_isvec; // @[LSU.scala 133:21]
  reg  reg_save_ctrl_mem_unsigned; // @[LSU.scala 133:21]
  reg [1:0] reg_save_ctrl_mem_cmd; // @[LSU.scala 133:21]
  reg [1:0] reg_save_ctrl_mop; // @[LSU.scala 133:21]
  reg [4:0] reg_save_ctrl_reg_idxw; // @[LSU.scala 133:21]
  reg  reg_save_ctrl_wfd; // @[LSU.scala 133:21]
  reg  reg_save_ctrl_wxd; // @[LSU.scala 133:21]
  reg [1:0] reg_entryID; // @[LSU.scala 136:28]
  wire [32:0] _addr_0_T_3 = 1'h0 * reg_save_in2_0; // @[LSU.scala 146:61]
  wire [32:0] _addr_0_T_4 = reg_save_ctrl_mop == 2'h3 ? {{1'd0}, reg_save_in2_0} : _addr_0_T_3; // @[LSU.scala 146:12]
  wire [32:0] _addr_0_T_5 = reg_save_ctrl_mop == 2'h0 ? 33'h0 : _addr_0_T_4; // @[LSU.scala 145:28]
  wire [32:0] _GEN_201 = {{1'd0}, reg_save_in1_0}; // @[LSU.scala 145:23]
  wire [32:0] _addr_0_T_7 = _GEN_201 + _addr_0_T_5; // @[LSU.scala 145:23]
  wire [31:0] _addr_0_T_9 = reg_save_in1_0 + reg_save_in2_0; // @[LSU.scala 147:23]
  wire [32:0] _addr_0_T_10 = reg_save_ctrl_isvec ? _addr_0_T_7 : {{1'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_0 = _addr_0_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_0 = ~reg_save_mask_0 | addr_0 < 32'h1000; // @[LSU.scala 149:39]
  wire [32:0] _addr_1_T_3 = 1'h1 * reg_save_in2_1; // @[LSU.scala 146:61]
  wire [32:0] _addr_1_T_4 = reg_save_ctrl_mop == 2'h3 ? {{1'd0}, reg_save_in2_1} : _addr_1_T_3; // @[LSU.scala 146:12]
  wire [32:0] _addr_1_T_5 = reg_save_ctrl_mop == 2'h0 ? 33'h4 : _addr_1_T_4; // @[LSU.scala 145:28]
  wire [32:0] _GEN_202 = {{1'd0}, reg_save_in1_1}; // @[LSU.scala 145:23]
  wire [32:0] _addr_1_T_7 = _GEN_202 + _addr_1_T_5; // @[LSU.scala 145:23]
  wire [32:0] _addr_1_T_10 = reg_save_ctrl_isvec ? _addr_1_T_7 : {{1'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_1 = _addr_1_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_1 = ~reg_save_mask_1 | addr_1 < 32'h1000; // @[LSU.scala 149:39]
  wire [33:0] _addr_2_T_3 = 2'h2 * reg_save_in2_2; // @[LSU.scala 146:61]
  wire [33:0] _addr_2_T_4 = reg_save_ctrl_mop == 2'h3 ? {{2'd0}, reg_save_in2_2} : _addr_2_T_3; // @[LSU.scala 146:12]
  wire [33:0] _addr_2_T_5 = reg_save_ctrl_mop == 2'h0 ? 34'h8 : _addr_2_T_4; // @[LSU.scala 145:28]
  wire [33:0] _GEN_203 = {{2'd0}, reg_save_in1_2}; // @[LSU.scala 145:23]
  wire [33:0] _addr_2_T_7 = _GEN_203 + _addr_2_T_5; // @[LSU.scala 145:23]
  wire [33:0] _addr_2_T_10 = reg_save_ctrl_isvec ? _addr_2_T_7 : {{2'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_2 = _addr_2_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_2 = ~reg_save_mask_2 | addr_2 < 32'h1000; // @[LSU.scala 149:39]
  wire [33:0] _addr_3_T_3 = 2'h3 * reg_save_in2_3; // @[LSU.scala 146:61]
  wire [33:0] _addr_3_T_4 = reg_save_ctrl_mop == 2'h3 ? {{2'd0}, reg_save_in2_3} : _addr_3_T_3; // @[LSU.scala 146:12]
  wire [33:0] _addr_3_T_5 = reg_save_ctrl_mop == 2'h0 ? 34'hc : _addr_3_T_4; // @[LSU.scala 145:28]
  wire [33:0] _GEN_204 = {{2'd0}, reg_save_in1_3}; // @[LSU.scala 145:23]
  wire [33:0] _addr_3_T_7 = _GEN_204 + _addr_3_T_5; // @[LSU.scala 145:23]
  wire [33:0] _addr_3_T_10 = reg_save_ctrl_isvec ? _addr_3_T_7 : {{2'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_3 = _addr_3_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_3 = ~reg_save_mask_3 | addr_3 < 32'h1000; // @[LSU.scala 149:39]
  wire [34:0] _addr_4_T_3 = 3'h4 * reg_save_in2_4; // @[LSU.scala 146:61]
  wire [34:0] _addr_4_T_4 = reg_save_ctrl_mop == 2'h3 ? {{3'd0}, reg_save_in2_4} : _addr_4_T_3; // @[LSU.scala 146:12]
  wire [34:0] _addr_4_T_5 = reg_save_ctrl_mop == 2'h0 ? 35'h10 : _addr_4_T_4; // @[LSU.scala 145:28]
  wire [34:0] _GEN_205 = {{3'd0}, reg_save_in1_4}; // @[LSU.scala 145:23]
  wire [34:0] _addr_4_T_7 = _GEN_205 + _addr_4_T_5; // @[LSU.scala 145:23]
  wire [34:0] _addr_4_T_10 = reg_save_ctrl_isvec ? _addr_4_T_7 : {{3'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_4 = _addr_4_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_4 = ~reg_save_mask_4 | addr_4 < 32'h1000; // @[LSU.scala 149:39]
  wire [34:0] _addr_5_T_3 = 3'h5 * reg_save_in2_5; // @[LSU.scala 146:61]
  wire [34:0] _addr_5_T_4 = reg_save_ctrl_mop == 2'h3 ? {{3'd0}, reg_save_in2_5} : _addr_5_T_3; // @[LSU.scala 146:12]
  wire [34:0] _addr_5_T_5 = reg_save_ctrl_mop == 2'h0 ? 35'h14 : _addr_5_T_4; // @[LSU.scala 145:28]
  wire [34:0] _GEN_206 = {{3'd0}, reg_save_in1_5}; // @[LSU.scala 145:23]
  wire [34:0] _addr_5_T_7 = _GEN_206 + _addr_5_T_5; // @[LSU.scala 145:23]
  wire [34:0] _addr_5_T_10 = reg_save_ctrl_isvec ? _addr_5_T_7 : {{3'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_5 = _addr_5_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_5 = ~reg_save_mask_5 | addr_5 < 32'h1000; // @[LSU.scala 149:39]
  wire [34:0] _addr_6_T_3 = 3'h6 * reg_save_in2_6; // @[LSU.scala 146:61]
  wire [34:0] _addr_6_T_4 = reg_save_ctrl_mop == 2'h3 ? {{3'd0}, reg_save_in2_6} : _addr_6_T_3; // @[LSU.scala 146:12]
  wire [34:0] _addr_6_T_5 = reg_save_ctrl_mop == 2'h0 ? 35'h18 : _addr_6_T_4; // @[LSU.scala 145:28]
  wire [34:0] _GEN_207 = {{3'd0}, reg_save_in1_6}; // @[LSU.scala 145:23]
  wire [34:0] _addr_6_T_7 = _GEN_207 + _addr_6_T_5; // @[LSU.scala 145:23]
  wire [34:0] _addr_6_T_10 = reg_save_ctrl_isvec ? _addr_6_T_7 : {{3'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_6 = _addr_6_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_6 = ~reg_save_mask_6 | addr_6 < 32'h1000; // @[LSU.scala 149:39]
  wire [34:0] _addr_7_T_3 = 3'h7 * reg_save_in2_7; // @[LSU.scala 146:61]
  wire [34:0] _addr_7_T_4 = reg_save_ctrl_mop == 2'h3 ? {{3'd0}, reg_save_in2_7} : _addr_7_T_3; // @[LSU.scala 146:12]
  wire [34:0] _addr_7_T_5 = reg_save_ctrl_mop == 2'h0 ? 35'h1c : _addr_7_T_4; // @[LSU.scala 145:28]
  wire [34:0] _GEN_208 = {{3'd0}, reg_save_in1_7}; // @[LSU.scala 145:23]
  wire [34:0] _addr_7_T_7 = _GEN_208 + _addr_7_T_5; // @[LSU.scala 145:23]
  wire [34:0] _addr_7_T_10 = reg_save_ctrl_isvec ? _addr_7_T_7 : {{3'd0}, _addr_0_T_9}; // @[LSU.scala 144:19]
  wire [31:0] addr_7 = _addr_7_T_10[31:0]; // @[LSU.scala 138:18 144:13]
  wire  is_shared_7 = ~reg_save_mask_7 | addr_7 < 32'h1000; // @[LSU.scala 149:39]
  wire [7:0] _all_shared_T = {is_shared_7,is_shared_6,is_shared_5,is_shared_4,is_shared_3,is_shared_2,is_shared_1,
    is_shared_0}; // @[LSU.scala 152:15]
  wire  _all_shared_T_1 = &_all_shared_T; // @[LSU.scala 152:22]
  wire  all_shared = reg_save_ctrl_isvec ? _all_shared_T_1 : is_shared_0; // @[LSU.scala 151:20]
  wire [7:0] _addr_wire_T = {reg_save_mask_7,reg_save_mask_6,reg_save_mask_5,reg_save_mask_4,reg_save_mask_3,
    reg_save_mask_2,reg_save_mask_1,reg_save_mask_0}; // @[LSU.scala 156:49]
  wire [2:0] _addr_wire_T_9 = _addr_wire_T[6] ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _addr_wire_T_10 = _addr_wire_T[5] ? 3'h5 : _addr_wire_T_9; // @[Mux.scala 47:70]
  wire [2:0] _addr_wire_T_11 = _addr_wire_T[4] ? 3'h4 : _addr_wire_T_10; // @[Mux.scala 47:70]
  wire [2:0] _addr_wire_T_12 = _addr_wire_T[3] ? 3'h3 : _addr_wire_T_11; // @[Mux.scala 47:70]
  wire [2:0] _addr_wire_T_13 = _addr_wire_T[2] ? 3'h2 : _addr_wire_T_12; // @[Mux.scala 47:70]
  wire [2:0] _addr_wire_T_14 = _addr_wire_T[1] ? 3'h1 : _addr_wire_T_13; // @[Mux.scala 47:70]
  wire [2:0] _addr_wire_T_15 = _addr_wire_T[0] ? 3'h0 : _addr_wire_T_14; // @[Mux.scala 47:70]
  wire [31:0] _GEN_1 = 3'h1 == _addr_wire_T_15 ? addr_1 : addr_0; // @[LSU.scala 156:{12,12}]
  wire [31:0] _GEN_2 = 3'h2 == _addr_wire_T_15 ? addr_2 : _GEN_1; // @[LSU.scala 156:{12,12}]
  wire [31:0] _GEN_3 = 3'h3 == _addr_wire_T_15 ? addr_3 : _GEN_2; // @[LSU.scala 156:{12,12}]
  wire [31:0] _GEN_4 = 3'h4 == _addr_wire_T_15 ? addr_4 : _GEN_3; // @[LSU.scala 156:{12,12}]
  wire [31:0] _GEN_5 = 3'h5 == _addr_wire_T_15 ? addr_5 : _GEN_4; // @[LSU.scala 156:{12,12}]
  wire [31:0] _GEN_6 = 3'h6 == _addr_wire_T_15 ? addr_6 : _GEN_5; // @[LSU.scala 156:{12,12}]
  wire [31:0] addr_wire = 3'h7 == _addr_wire_T_15 ? addr_7 : _GEN_6; // @[LSU.scala 156:{12,12}]
  wire  _tag_T_1 = _addr_wire_T != 8'h0; // @[LSU.scala 157:39]
  wire [21:0] tag = _addr_wire_T != 8'h0 ? addr_wire[31:10] : 22'h0; // @[LSU.scala 157:16]
  wire [4:0] setIdx = _tag_T_1 ? addr_wire[9:5] : 5'h0; // @[LSU.scala 158:19]
  wire  _io_to_mshr_valid_T_1 = |reg_save_ctrl_mem_cmd; // @[LSU.scala 190:63]
  wire  _io_to_shared_bits_perLaneAddr_0_activeMask_T_4 = addr_0[31:10] == tag & addr_0[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_1_activeMask_T_4 = addr_1[31:10] == tag & addr_1[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_2_activeMask_T_4 = addr_2[31:10] == tag & addr_2[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_3_activeMask_T_4 = addr_3[31:10] == tag & addr_3[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_4_activeMask_T_4 = addr_4[31:10] == tag & addr_4[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_5_activeMask_T_4 = addr_5[31:10] == tag & addr_5[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_6_activeMask_T_4 = addr_6[31:10] == tag & addr_6[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  _io_to_shared_bits_perLaneAddr_7_activeMask_T_4 = addr_7[31:10] == tag & addr_7[9:5] == setIdx; // @[LSU.scala 203:120]
  wire  mask_next_0 = reg_save_mask_0 & ~_io_to_shared_bits_perLaneAddr_0_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_1 = reg_save_mask_1 & ~_io_to_shared_bits_perLaneAddr_1_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_2 = reg_save_mask_2 & ~_io_to_shared_bits_perLaneAddr_2_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_3 = reg_save_mask_3 & ~_io_to_shared_bits_perLaneAddr_3_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_4 = reg_save_mask_4 & ~_io_to_shared_bits_perLaneAddr_4_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_5 = reg_save_mask_5 & ~_io_to_shared_bits_perLaneAddr_5_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_6 = reg_save_mask_6 & ~_io_to_shared_bits_perLaneAddr_6_activeMask_T_4; // @[LSU.scala 224:38]
  wire  mask_next_7 = reg_save_mask_7 & ~_io_to_shared_bits_perLaneAddr_7_activeMask_T_4; // @[LSU.scala 224:38]
  wire  _T_24 = 2'h0 == state; // @[LSU.scala 229:16]
  wire  _T_25 = 2'h1 == state; // @[LSU.scala 229:16]
  wire  _T_27 = io_to_mshr_ready & io_to_mshr_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_9 = _T_27 ? 2'h2 : 2'h1; // @[LSU.scala 237:{34,41,70}]
  wire [1:0] _GEN_10 = _T_27 ? 2'h3 : 2'h1; // @[LSU.scala 239:{34,41,70}]
  wire [1:0] _GEN_11 = all_shared ? _GEN_9 : _GEN_10; // @[LSU.scala 236:25]
  wire  _T_29 = 2'h2 == state; // @[LSU.scala 229:16]
  wire  _T_30 = io_to_shared_ready & io_to_shared_valid; // @[Decoupled.scala 50:35]
  wire [7:0] _T_32 = {mask_next_7,mask_next_6,mask_next_5,mask_next_4,mask_next_3,mask_next_2,mask_next_1,mask_next_0}; // @[LSU.scala 245:57]
  wire  _T_33 = _T_32 == 8'h0; // @[LSU.scala 245:59]
  wire [1:0] _GEN_14 = _T_32 == 8'h0 ? 2'h0 : 2'h2; // @[LSU.scala 245:66 246:30 248:28]
  wire [1:0] _GEN_16 = _T_30 ? _GEN_14 : 2'h2; // @[LSU.scala 244:32 250:25]
  wire  _T_35 = 2'h3 == state; // @[LSU.scala 229:16]
  wire  _T_36 = io_to_dcache_ready & io_to_dcache_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_18 = _T_33 ? 2'h0 : 2'h3; // @[LSU.scala 254:66 255:30 257:28]
  wire [1:0] _GEN_20 = _T_36 ? _GEN_18 : 2'h3; // @[LSU.scala 253:32 259:25]
  wire [1:0] _GEN_22 = 2'h3 == state ? _GEN_20 : state; // @[LSU.scala 229:16 131:22]
  wire  _T_42 = io_from_fifo_ready & io_from_fifo_valid; // @[Decoupled.scala 50:35]
  wire  _T_43_0 = io_from_fifo_bits_ctrl_isvec ? io_from_fifo_bits_mask_0 : 1'h1; // @[LSU.scala 267:29]
  wire  _GEN_30 = _T_42 & io_from_fifo_bits_ctrl_wxd; // @[LSU.scala 265:32 266:18 268:28]
  wire  _GEN_35 = _T_42 & io_from_fifo_bits_ctrl_wfd; // @[LSU.scala 265:32 266:18 268:28]
  wire  _GEN_44 = _T_42 & io_from_fifo_bits_ctrl_mem_unsigned; // @[LSU.scala 265:32 266:18 268:28]
  wire  _GEN_49 = _T_42 & io_from_fifo_bits_ctrl_isvec; // @[LSU.scala 265:32 266:18 268:28]
  wire  _GEN_61 = _T_42 & _T_43_0; // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_62 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_1); // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_63 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_2); // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_64 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_3); // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_65 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_4); // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_66 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_5); // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_67 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_6); // @[LSU.scala 265:32 267:23 268:28]
  wire  _GEN_68 = _T_42 & (io_from_fifo_bits_ctrl_isvec & io_from_fifo_bits_mask_7); // @[LSU.scala 265:32 267:23 268:28]
  wire [1:0] _GEN_93 = _T_27 ? io_idx_entry : reg_entryID; // @[LSU.scala 136:28 272:{32,45}]
  wire  _GEN_103 = _T_36 ? mask_next_0 : reg_save_mask_0; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_104 = _T_36 ? mask_next_1 : reg_save_mask_1; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_105 = _T_36 ? mask_next_2 : reg_save_mask_2; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_106 = _T_36 ? mask_next_3 : reg_save_mask_3; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_107 = _T_36 ? mask_next_4 : reg_save_mask_4; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_108 = _T_36 ? mask_next_5 : reg_save_mask_5; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_109 = _T_36 ? mask_next_6 : reg_save_mask_6; // @[LSU.scala 284:32 285:23 287:23]
  wire  _GEN_110 = _T_36 ? mask_next_7 : reg_save_mask_7; // @[LSU.scala 284:32 285:23 287:23]
  assign io_from_fifo_ready = state == 2'h0; // @[LSU.scala 135:30]
  assign io_to_mshr_valid = state == 2'h1 & |reg_save_ctrl_mem_cmd; // @[LSU.scala 190:38]
  assign io_to_mshr_bits_tag_warp_id = reg_save_ctrl_wid; // @[LSU.scala 184:31]
  assign io_to_mshr_bits_tag_wfd = reg_save_ctrl_wfd; // @[LSU.scala 186:26]
  assign io_to_mshr_bits_tag_wxd = reg_save_ctrl_wxd; // @[LSU.scala 185:26]
  assign io_to_mshr_bits_tag_reg_idxw = reg_save_ctrl_reg_idxw; // @[LSU.scala 183:32]
  assign io_to_mshr_bits_tag_mask_0 = reg_save_mask_0; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_1 = reg_save_mask_1; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_2 = reg_save_mask_2; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_3 = reg_save_mask_3; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_4 = reg_save_mask_4; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_5 = reg_save_mask_5; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_6 = reg_save_mask_6; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_mask_7 = reg_save_mask_7; // @[LSU.scala 182:28]
  assign io_to_mshr_bits_tag_unsigned = reg_save_ctrl_mem_unsigned; // @[LSU.scala 188:32]
  assign io_to_mshr_bits_tag_isvec = reg_save_ctrl_isvec; // @[LSU.scala 187:29]
  assign io_to_mshr_bits_tag_isWrite = reg_save_ctrl_mem_cmd[1]; // @[LSU.scala 191:55]
  assign io_to_dcache_valid = state == 2'h3; // @[LSU.scala 221:30]
  assign io_to_dcache_bits_instrId = reg_entryID; // @[LSU.scala 210:29]
  assign io_to_dcache_bits_isWrite = reg_save_ctrl_mem_cmd[1]; // @[LSU.scala 220:53]
  assign io_to_dcache_bits_tag = _addr_wire_T != 8'h0 ? addr_wire[31:10] : 22'h0; // @[LSU.scala 157:16]
  assign io_to_dcache_bits_setIdx = _tag_T_1 ? addr_wire[9:5] : 5'h0; // @[LSU.scala 158:19]
  assign io_to_dcache_bits_perLaneAddr_0_activeMask = reg_save_mask_0 & _io_to_shared_bits_perLaneAddr_0_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_0_blockOffset = addr_0[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_1_activeMask = reg_save_mask_1 & _io_to_shared_bits_perLaneAddr_1_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_1_blockOffset = addr_1[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_2_activeMask = reg_save_mask_2 & _io_to_shared_bits_perLaneAddr_2_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_2_blockOffset = addr_2[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_3_activeMask = reg_save_mask_3 & _io_to_shared_bits_perLaneAddr_3_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_3_blockOffset = addr_3[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_4_activeMask = reg_save_mask_4 & _io_to_shared_bits_perLaneAddr_4_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_4_blockOffset = addr_4[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_5_activeMask = reg_save_mask_5 & _io_to_shared_bits_perLaneAddr_5_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_5_blockOffset = addr_5[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_6_activeMask = reg_save_mask_6 & _io_to_shared_bits_perLaneAddr_6_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_6_blockOffset = addr_6[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_perLaneAddr_7_activeMask = reg_save_mask_7 & _io_to_shared_bits_perLaneAddr_7_activeMask_T_4; // @[LSU.scala 217:69]
  assign io_to_dcache_bits_perLaneAddr_7_blockOffset = addr_7[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_dcache_bits_data_0 = reg_save_in3_0; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_1 = reg_save_in3_1; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_2 = reg_save_in3_2; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_3 = reg_save_in3_3; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_4 = reg_save_in3_4; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_5 = reg_save_in3_5; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_6 = reg_save_in3_6; // @[LSU.scala 219:26]
  assign io_to_dcache_bits_data_7 = reg_save_in3_7; // @[LSU.scala 219:26]
  assign io_to_shared_valid = state == 2'h2; // @[LSU.scala 207:30]
  assign io_to_shared_bits_instrId = reg_entryID; // @[LSU.scala 196:29]
  assign io_to_shared_bits_isWrite = reg_save_ctrl_mem_cmd[1]; // @[LSU.scala 206:53]
  assign io_to_shared_bits_setIdx = _tag_T_1 ? addr_wire[9:5] : 5'h0; // @[LSU.scala 158:19]
  assign io_to_shared_bits_perLaneAddr_0_activeMask = reg_save_mask_0 & (addr_0[31:10] == tag & addr_0[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_0_blockOffset = addr_0[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_1_activeMask = reg_save_mask_1 & (addr_1[31:10] == tag & addr_1[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_1_blockOffset = addr_1[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_2_activeMask = reg_save_mask_2 & (addr_2[31:10] == tag & addr_2[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_2_blockOffset = addr_2[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_3_activeMask = reg_save_mask_3 & (addr_3[31:10] == tag & addr_3[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_3_blockOffset = addr_3[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_4_activeMask = reg_save_mask_4 & (addr_4[31:10] == tag & addr_4[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_4_blockOffset = addr_4[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_5_activeMask = reg_save_mask_5 & (addr_5[31:10] == tag & addr_5[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_5_blockOffset = addr_5[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_6_activeMask = reg_save_mask_6 & (addr_6[31:10] == tag & addr_6[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_6_blockOffset = addr_6[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_perLaneAddr_7_activeMask = reg_save_mask_7 & (addr_7[31:10] == tag & addr_7[9:5] == setIdx); // @[LSU.scala 203:69]
  assign io_to_shared_bits_perLaneAddr_7_blockOffset = addr_7[4:2]; // @[LSU.scala 163:25 164:55]
  assign io_to_shared_bits_data_0 = reg_save_in3_0; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_1 = reg_save_in3_1; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_2 = reg_save_in3_2; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_3 = reg_save_in3_3; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_4 = reg_save_in3_4; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_5 = reg_save_in3_5; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_6 = reg_save_in3_6; // @[LSU.scala 205:26]
  assign io_to_shared_bits_data_7 = reg_save_in3_7; // @[LSU.scala 205:26]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 131:22]
      state <= 2'h0; // @[LSU.scala 131:22]
    end else if (2'h0 == state) begin // @[LSU.scala 229:16]
      if (io_from_fifo_valid) begin // @[LSU.scala 231:31]
        state <= 2'h1; // @[LSU.scala 231:39]
      end
    end else if (2'h1 == state) begin // @[LSU.scala 229:16]
      if (_io_to_mshr_valid_T_1) begin // @[LSU.scala 235:38]
        state <= _GEN_11;
      end else begin
        state <= 2'h0; // @[LSU.scala 241:26]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 229:16]
      state <= _GEN_16;
    end else begin
      state <= _GEN_22;
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_0 <= io_from_fifo_bits_in1_0; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_0 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_1 <= io_from_fifo_bits_in1_1; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_1 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_2 <= io_from_fifo_bits_in1_2; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_2 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_3 <= io_from_fifo_bits_in1_3; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_3 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_4 <= io_from_fifo_bits_in1_4; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_4 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_5 <= io_from_fifo_bits_in1_5; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_5 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_6 <= io_from_fifo_bits_in1_6; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_6 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in1_7 <= io_from_fifo_bits_in1_7; // @[LSU.scala 266:18]
      end else begin
        reg_save_in1_7 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_0 <= io_from_fifo_bits_in2_0; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_0 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_1 <= io_from_fifo_bits_in2_1; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_1 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_2 <= io_from_fifo_bits_in2_2; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_2 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_3 <= io_from_fifo_bits_in2_3; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_3 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_4 <= io_from_fifo_bits_in2_4; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_4 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_5 <= io_from_fifo_bits_in2_5; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_5 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_6 <= io_from_fifo_bits_in2_6; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_6 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in2_7 <= io_from_fifo_bits_in2_7; // @[LSU.scala 266:18]
      end else begin
        reg_save_in2_7 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_0 <= io_from_fifo_bits_in3_0; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_0 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_1 <= io_from_fifo_bits_in3_1; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_1 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_2 <= io_from_fifo_bits_in3_2; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_2 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_3 <= io_from_fifo_bits_in3_3; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_3 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_4 <= io_from_fifo_bits_in3_4; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_4 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_5 <= io_from_fifo_bits_in3_5; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_5 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_6 <= io_from_fifo_bits_in3_6; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_6 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_in3_7 <= io_from_fifo_bits_in3_7; // @[LSU.scala 266:18]
      end else begin
        reg_save_in3_7 <= 32'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_0 <= _GEN_61;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_0 <= mask_next_0; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_0 <= _GEN_103;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_1 <= _GEN_62;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_1 <= mask_next_1; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_1 <= _GEN_104;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_2 <= _GEN_63;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_2 <= mask_next_2; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_2 <= _GEN_105;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_3 <= _GEN_64;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_3 <= mask_next_3; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_3 <= _GEN_106;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_4 <= _GEN_65;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_4 <= mask_next_4; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_4 <= _GEN_107;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_5 <= _GEN_66;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_5 <= mask_next_5; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_5 <= _GEN_108;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_6 <= _GEN_67;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_6 <= mask_next_6; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_6 <= _GEN_109;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_mask_7 <= _GEN_68;
    end else if (!(_T_25)) begin // @[LSU.scala 263:16]
      if (_T_29) begin // @[LSU.scala 263:16]
        if (_T_30) begin // @[LSU.scala 277:32]
          reg_save_mask_7 <= mask_next_7; // @[LSU.scala 278:23]
        end
      end else if (_T_35) begin // @[LSU.scala 263:16]
        reg_save_mask_7 <= _GEN_110;
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_ctrl_wid <= io_from_fifo_bits_ctrl_wid; // @[LSU.scala 266:18]
      end else begin
        reg_save_ctrl_wid <= 2'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_ctrl_isvec <= _GEN_49;
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_ctrl_mem_unsigned <= _GEN_44;
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_ctrl_mem_cmd <= io_from_fifo_bits_ctrl_mem_cmd; // @[LSU.scala 266:18]
      end else begin
        reg_save_ctrl_mem_cmd <= 2'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_ctrl_mop <= io_from_fifo_bits_ctrl_mop; // @[LSU.scala 266:18]
      end else begin
        reg_save_ctrl_mop <= 2'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      if (_T_42) begin // @[LSU.scala 265:32]
        reg_save_ctrl_reg_idxw <= io_from_fifo_bits_ctrl_reg_idxw; // @[LSU.scala 266:18]
      end else begin
        reg_save_ctrl_reg_idxw <= 5'h0; // @[LSU.scala 268:28]
      end
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_ctrl_wfd <= _GEN_35;
    end
    if (_T_24) begin // @[LSU.scala 263:16]
      reg_save_ctrl_wxd <= _GEN_30;
    end
    if (reset) begin // @[LSU.scala 136:28]
      reg_entryID <= 2'h0; // @[LSU.scala 136:28]
    end else if (!(_T_24)) begin // @[LSU.scala 263:16]
      if (_T_25) begin // @[LSU.scala 263:16]
        if (_io_to_mshr_valid_T_1) begin // @[LSU.scala 271:38]
          reg_entryID <= _GEN_93;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reg_save_in1_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_save_in1_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_save_in1_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_save_in1_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_save_in1_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_save_in1_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_save_in1_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_save_in1_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_save_in2_0 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_save_in2_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_save_in2_2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_save_in2_3 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_save_in2_4 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_save_in2_5 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_save_in2_6 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_save_in2_7 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_save_in3_0 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_save_in3_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_save_in3_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_save_in3_3 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_save_in3_4 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_save_in3_5 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_save_in3_6 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_save_in3_7 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_save_mask_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  reg_save_mask_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  reg_save_mask_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  reg_save_mask_3 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  reg_save_mask_4 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  reg_save_mask_5 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  reg_save_mask_6 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  reg_save_mask_7 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  reg_save_ctrl_wid = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  reg_save_ctrl_isvec = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  reg_save_ctrl_mem_unsigned = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  reg_save_ctrl_mem_cmd = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  reg_save_ctrl_mop = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  reg_save_ctrl_reg_idxw = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  reg_save_ctrl_wfd = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  reg_save_ctrl_wxd = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  reg_entryID = _RAND_41[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_8(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_instrId,
  input  [31:0] io_in_0_bits_data_0,
  input  [31:0] io_in_0_bits_data_1,
  input  [31:0] io_in_0_bits_data_2,
  input  [31:0] io_in_0_bits_data_3,
  input  [31:0] io_in_0_bits_data_4,
  input  [31:0] io_in_0_bits_data_5,
  input  [31:0] io_in_0_bits_data_6,
  input  [31:0] io_in_0_bits_data_7,
  input         io_in_0_bits_activeMask_0,
  input         io_in_0_bits_activeMask_1,
  input         io_in_0_bits_activeMask_2,
  input         io_in_0_bits_activeMask_3,
  input         io_in_0_bits_activeMask_4,
  input         io_in_0_bits_activeMask_5,
  input         io_in_0_bits_activeMask_6,
  input         io_in_0_bits_activeMask_7,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_instrId,
  input  [31:0] io_in_1_bits_data_0,
  input  [31:0] io_in_1_bits_data_1,
  input  [31:0] io_in_1_bits_data_2,
  input  [31:0] io_in_1_bits_data_3,
  input  [31:0] io_in_1_bits_data_4,
  input  [31:0] io_in_1_bits_data_5,
  input  [31:0] io_in_1_bits_data_6,
  input  [31:0] io_in_1_bits_data_7,
  input         io_in_1_bits_activeMask_0,
  input         io_in_1_bits_activeMask_1,
  input         io_in_1_bits_activeMask_2,
  input         io_in_1_bits_activeMask_3,
  input         io_in_1_bits_activeMask_4,
  input         io_in_1_bits_activeMask_5,
  input         io_in_1_bits_activeMask_6,
  input         io_in_1_bits_activeMask_7,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_instrId,
  output [31:0] io_out_bits_data_0,
  output [31:0] io_out_bits_data_1,
  output [31:0] io_out_bits_data_2,
  output [31:0] io_out_bits_data_3,
  output [31:0] io_out_bits_data_4,
  output [31:0] io_out_bits_data_5,
  output [31:0] io_out_bits_data_6,
  output [31:0] io_out_bits_data_7,
  output        io_out_bits_activeMask_0,
  output        io_out_bits_activeMask_1,
  output        io_out_bits_activeMask_2,
  output        io_out_bits_activeMask_3,
  output        io_out_bits_activeMask_4,
  output        io_out_bits_activeMask_5,
  output        io_out_bits_activeMask_6,
  output        io_out_bits_activeMask_7
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_instrId = io_in_0_valid ? io_in_0_bits_instrId : io_in_1_bits_instrId; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_0 = io_in_0_valid ? io_in_0_bits_data_0 : io_in_1_bits_data_0; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_1 = io_in_0_valid ? io_in_0_bits_data_1 : io_in_1_bits_data_1; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_2 = io_in_0_valid ? io_in_0_bits_data_2 : io_in_1_bits_data_2; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_3 = io_in_0_valid ? io_in_0_bits_data_3 : io_in_1_bits_data_3; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_4 = io_in_0_valid ? io_in_0_bits_data_4 : io_in_1_bits_data_4; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_5 = io_in_0_valid ? io_in_0_bits_data_5 : io_in_1_bits_data_5; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_6 = io_in_0_valid ? io_in_0_bits_data_6 : io_in_1_bits_data_6; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data_7 = io_in_0_valid ? io_in_0_bits_data_7 : io_in_1_bits_data_7; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_0 = io_in_0_valid ? io_in_0_bits_activeMask_0 : io_in_1_bits_activeMask_0; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_1 = io_in_0_valid ? io_in_0_bits_activeMask_1 : io_in_1_bits_activeMask_1; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_2 = io_in_0_valid ? io_in_0_bits_activeMask_2 : io_in_1_bits_activeMask_2; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_3 = io_in_0_valid ? io_in_0_bits_activeMask_3 : io_in_1_bits_activeMask_3; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_4 = io_in_0_valid ? io_in_0_bits_activeMask_4 : io_in_1_bits_activeMask_4; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_5 = io_in_0_valid ? io_in_0_bits_activeMask_5 : io_in_1_bits_activeMask_5; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_6 = io_in_0_valid ? io_in_0_bits_activeMask_6 : io_in_1_bits_activeMask_6; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_activeMask_7 = io_in_0_valid ? io_in_0_bits_activeMask_7 : io_in_1_bits_activeMask_7; // @[Arbiter.scala 139:15 141:26 143:19]
endmodule
module MSHRv2(
  input         clock,
  input         reset,
  output        io_from_addr_ready,
  input         io_from_addr_valid,
  input  [1:0]  io_from_addr_bits_tag_warp_id,
  input         io_from_addr_bits_tag_wfd,
  input         io_from_addr_bits_tag_wxd,
  input  [4:0]  io_from_addr_bits_tag_reg_idxw,
  input         io_from_addr_bits_tag_mask_0,
  input         io_from_addr_bits_tag_mask_1,
  input         io_from_addr_bits_tag_mask_2,
  input         io_from_addr_bits_tag_mask_3,
  input         io_from_addr_bits_tag_mask_4,
  input         io_from_addr_bits_tag_mask_5,
  input         io_from_addr_bits_tag_mask_6,
  input         io_from_addr_bits_tag_mask_7,
  input         io_from_addr_bits_tag_unsigned,
  input         io_from_addr_bits_tag_isvec,
  input         io_from_addr_bits_tag_isWrite,
  output [1:0]  io_idx_entry,
  output        io_from_dcache_ready,
  input         io_from_dcache_valid,
  input  [1:0]  io_from_dcache_bits_instrId,
  input  [31:0] io_from_dcache_bits_data_0,
  input  [31:0] io_from_dcache_bits_data_1,
  input  [31:0] io_from_dcache_bits_data_2,
  input  [31:0] io_from_dcache_bits_data_3,
  input  [31:0] io_from_dcache_bits_data_4,
  input  [31:0] io_from_dcache_bits_data_5,
  input  [31:0] io_from_dcache_bits_data_6,
  input  [31:0] io_from_dcache_bits_data_7,
  input         io_from_dcache_bits_activeMask_0,
  input         io_from_dcache_bits_activeMask_1,
  input         io_from_dcache_bits_activeMask_2,
  input         io_from_dcache_bits_activeMask_3,
  input         io_from_dcache_bits_activeMask_4,
  input         io_from_dcache_bits_activeMask_5,
  input         io_from_dcache_bits_activeMask_6,
  input         io_from_dcache_bits_activeMask_7,
  input         io_to_pipe_ready,
  output        io_to_pipe_valid,
  output [1:0]  io_to_pipe_bits_tag_warp_id,
  output        io_to_pipe_bits_tag_wfd,
  output        io_to_pipe_bits_tag_wxd,
  output [4:0]  io_to_pipe_bits_tag_reg_idxw,
  output        io_to_pipe_bits_tag_mask_0,
  output        io_to_pipe_bits_tag_mask_1,
  output        io_to_pipe_bits_tag_mask_2,
  output        io_to_pipe_bits_tag_mask_3,
  output        io_to_pipe_bits_tag_mask_4,
  output        io_to_pipe_bits_tag_mask_5,
  output        io_to_pipe_bits_tag_mask_6,
  output        io_to_pipe_bits_tag_mask_7,
  output        io_to_pipe_bits_tag_isWrite,
  output [31:0] io_to_pipe_bits_data_0,
  output [31:0] io_to_pipe_bits_data_1,
  output [31:0] io_to_pipe_bits_data_2,
  output [31:0] io_to_pipe_bits_data_3,
  output [31:0] io_to_pipe_bits_data_4,
  output [31:0] io_to_pipe_bits_data_5,
  output [31:0] io_to_pipe_bits_data_6,
  output [31:0] io_to_pipe_bits_data_7
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_0 [0:3]; // @[MSHR.scala 21:17]
  wire  data_0_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_0_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_0_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_0_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_0_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_0_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_0_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_0_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_0_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_0_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_0_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_0_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_0_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_0_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_0_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_1 [0:3]; // @[MSHR.scala 21:17]
  wire  data_1_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_1_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_1_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_1_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_1_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_1_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_1_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_1_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_1_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_1_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_1_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_1_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_1_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_1_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_1_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_2 [0:3]; // @[MSHR.scala 21:17]
  wire  data_2_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_2_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_2_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_2_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_2_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_2_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_2_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_2_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_2_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_2_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_2_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_2_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_2_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_2_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_2_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_3 [0:3]; // @[MSHR.scala 21:17]
  wire  data_3_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_3_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_3_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_3_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_3_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_3_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_3_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_3_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_3_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_3_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_3_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_3_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_3_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_3_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_3_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_4 [0:3]; // @[MSHR.scala 21:17]
  wire  data_4_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_4_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_4_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_4_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_4_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_4_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_4_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_4_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_4_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_4_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_4_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_4_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_4_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_4_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_4_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_5 [0:3]; // @[MSHR.scala 21:17]
  wire  data_5_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_5_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_5_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_5_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_5_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_5_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_5_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_5_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_5_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_5_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_5_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_5_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_5_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_5_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_5_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_6 [0:3]; // @[MSHR.scala 21:17]
  wire  data_6_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_6_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_6_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_6_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_6_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_6_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_6_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_6_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_6_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_6_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_6_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_6_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_6_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_6_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_6_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [31:0] data_7 [0:3]; // @[MSHR.scala 21:17]
  wire  data_7_raw_data_en; // @[MSHR.scala 21:17]
  wire [1:0] data_7_raw_data_addr; // @[MSHR.scala 21:17]
  wire [31:0] data_7_raw_data_data; // @[MSHR.scala 21:17]
  wire [31:0] data_7_MPORT_data; // @[MSHR.scala 21:17]
  wire [1:0] data_7_MPORT_addr; // @[MSHR.scala 21:17]
  wire  data_7_MPORT_mask; // @[MSHR.scala 21:17]
  wire  data_7_MPORT_en; // @[MSHR.scala 21:17]
  wire [31:0] data_7_MPORT_2_data; // @[MSHR.scala 21:17]
  wire [1:0] data_7_MPORT_2_addr; // @[MSHR.scala 21:17]
  wire  data_7_MPORT_2_mask; // @[MSHR.scala 21:17]
  wire  data_7_MPORT_2_en; // @[MSHR.scala 21:17]
  wire [31:0] data_7_MPORT_4_data; // @[MSHR.scala 21:17]
  wire [1:0] data_7_MPORT_4_addr; // @[MSHR.scala 21:17]
  wire  data_7_MPORT_4_mask; // @[MSHR.scala 21:17]
  wire  data_7_MPORT_4_en; // @[MSHR.scala 21:17]
  reg [51:0] tag [0:3]; // @[MSHR.scala 22:16]
  wire  tag_output_tag_MPORT_en; // @[MSHR.scala 22:16]
  wire [1:0] tag_output_tag_MPORT_addr; // @[MSHR.scala 22:16]
  wire [51:0] tag_output_tag_MPORT_data; // @[MSHR.scala 22:16]
  wire [51:0] tag_MPORT_1_data; // @[MSHR.scala 22:16]
  wire [1:0] tag_MPORT_1_addr; // @[MSHR.scala 22:16]
  wire  tag_MPORT_1_mask; // @[MSHR.scala 22:16]
  wire  tag_MPORT_1_en; // @[MSHR.scala 22:16]
  wire [51:0] tag_MPORT_3_data; // @[MSHR.scala 22:16]
  wire [1:0] tag_MPORT_3_addr; // @[MSHR.scala 22:16]
  wire  tag_MPORT_3_mask; // @[MSHR.scala 22:16]
  wire  tag_MPORT_3_en; // @[MSHR.scala 22:16]
  reg [7:0] currentMask_0; // @[MSHR.scala 24:28]
  reg [7:0] currentMask_1; // @[MSHR.scala 24:28]
  reg [7:0] currentMask_2; // @[MSHR.scala 24:28]
  reg [7:0] currentMask_3; // @[MSHR.scala 24:28]
  wire  _inv_activeMask_T = ~io_from_dcache_bits_activeMask_0; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_1 = ~io_from_dcache_bits_activeMask_1; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_2 = ~io_from_dcache_bits_activeMask_2; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_3 = ~io_from_dcache_bits_activeMask_3; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_4 = ~io_from_dcache_bits_activeMask_4; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_5 = ~io_from_dcache_bits_activeMask_5; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_6 = ~io_from_dcache_bits_activeMask_6; // @[MSHR.scala 25:67]
  wire  _inv_activeMask_T_7 = ~io_from_dcache_bits_activeMask_7; // @[MSHR.scala 25:67]
  wire [7:0] inv_activeMask = {_inv_activeMask_T_7,_inv_activeMask_T_6,_inv_activeMask_T_5,_inv_activeMask_T_4,
    _inv_activeMask_T_3,_inv_activeMask_T_2,_inv_activeMask_T_1,_inv_activeMask_T}; // @[MSHR.scala 25:72]
  reg [3:0] used; // @[MSHR.scala 26:21]
  wire [3:0] _complete_T_4 = {currentMask_3 == 8'h0,currentMask_2 == 8'h0,currentMask_1 == 8'h0,currentMask_0 == 8'h0}; // @[MSHR.scala 27:52]
  wire [3:0] complete = _complete_T_4 & used; // @[MSHR.scala 27:59]
  wire  _output_entry_T = |complete; // @[MSHR.scala 28:35]
  wire [1:0] _output_entry_T_5 = complete[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _output_entry_T_6 = complete[1] ? 2'h1 : _output_entry_T_5; // @[Mux.scala 47:70]
  wire [1:0] _output_entry_T_7 = complete[0] ? 2'h0 : _output_entry_T_6; // @[Mux.scala 47:70]
  wire [1:0] output_entry = |complete ? _output_entry_T_7 : 2'h0; // @[MSHR.scala 28:25]
  wire  _valid_entry_T = &used; // @[MSHR.scala 29:30]
  wire [3:0] _valid_entry_T_1 = ~used; // @[MSHR.scala 29:57]
  wire [1:0] _valid_entry_T_6 = _valid_entry_T_1[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _valid_entry_T_7 = _valid_entry_T_1[1] ? 2'h1 : _valid_entry_T_6; // @[Mux.scala 47:70]
  wire [1:0] _valid_entry_T_8 = _valid_entry_T_1[0] ? 2'h0 : _valid_entry_T_7; // @[Mux.scala 47:70]
  wire [1:0] valid_entry = &used ? 2'h0 : _valid_entry_T_8; // @[MSHR.scala 29:24]
  reg  reg_req_mask_0; // @[MSHR.scala 30:20]
  reg  reg_req_mask_1; // @[MSHR.scala 30:20]
  reg  reg_req_mask_2; // @[MSHR.scala 30:20]
  reg  reg_req_mask_3; // @[MSHR.scala 30:20]
  reg  reg_req_mask_4; // @[MSHR.scala 30:20]
  reg  reg_req_mask_5; // @[MSHR.scala 30:20]
  reg  reg_req_mask_6; // @[MSHR.scala 30:20]
  reg  reg_req_mask_7; // @[MSHR.scala 30:20]
  reg [1:0] state; // @[MSHR.scala 33:22]
  wire  _io_from_dcache_ready_T = state == 2'h0; // @[MSHR.scala 35:32]
  wire  _io_idx_entry_T = io_from_addr_ready & io_from_addr_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = io_from_dcache_ready & io_from_dcache_valid; // @[Decoupled.scala 50:35]
  wire [7:0] _T_3 = {io_from_dcache_bits_activeMask_7,io_from_dcache_bits_activeMask_6,io_from_dcache_bits_activeMask_5,
    io_from_dcache_bits_activeMask_4,io_from_dcache_bits_activeMask_3,io_from_dcache_bits_activeMask_2,
    io_from_dcache_bits_activeMask_1,io_from_dcache_bits_activeMask_0}; // @[MSHR.scala 43:112]
  wire [7:0] _GEN_1 = 2'h1 == io_from_dcache_bits_instrId ? currentMask_1 : currentMask_0; // @[MSHR.scala 43:{78,78}]
  wire [7:0] _GEN_2 = 2'h2 == io_from_dcache_bits_instrId ? currentMask_2 : _GEN_1; // @[MSHR.scala 43:{78,78}]
  wire [7:0] _GEN_3 = 2'h3 == io_from_dcache_bits_instrId ? currentMask_3 : _GEN_2; // @[MSHR.scala 43:{78,78}]
  wire [1:0] _GEN_4 = io_to_pipe_ready & _GEN_3 == _T_3 ? 2'h2 : 2'h0; // @[MSHR.scala 43:119 44:15 45:25]
  wire  _T_8 = state == 2'h2; // @[MSHR.scala 51:19]
  wire [3:0] _T_9 = 4'h1 << valid_entry; // @[MSHR.scala 52:45]
  wire [3:0] _T_11 = ~complete; // @[MSHR.scala 52:45]
  wire [3:0] _T_12 = _T_11 | _T_9; // @[MSHR.scala 52:45]
  wire [3:0] _T_13 = ~_T_12; // @[MSHR.scala 52:45]
  wire [1:0] _GEN_9 = io_to_pipe_ready & _output_entry_T ? 2'h2 : 2'h0; // @[MSHR.scala 54:{43,49,73}]
  wire  _T_20 = 2'h0 == state; // @[MSHR.scala 57:16]
  wire [7:0] _currentMask_T = _GEN_3 & inv_activeMask; // @[MSHR.scala 61:94]
  wire [3:0] _used_T_1 = used | _T_9; // @[MSHR.scala 64:28]
  wire [34:0] lo_1 = {io_from_addr_bits_tag_unsigned,io_from_addr_bits_tag_isvec,4'hf,12'hfff,12'hfff,4'hf,
    io_from_addr_bits_tag_isWrite}; // @[MSHR.scala 67:33]
  wire [5:0] hi_lo_1 = {io_from_addr_bits_tag_mask_5,io_from_addr_bits_tag_mask_4,io_from_addr_bits_tag_mask_3,
    io_from_addr_bits_tag_mask_2,io_from_addr_bits_tag_mask_1,io_from_addr_bits_tag_mask_0}; // @[MSHR.scala 67:33]
  wire [16:0] hi_1 = {io_from_addr_bits_tag_warp_id,io_from_addr_bits_tag_wfd,io_from_addr_bits_tag_wxd,
    io_from_addr_bits_tag_reg_idxw,io_from_addr_bits_tag_mask_7,io_from_addr_bits_tag_mask_6,hi_lo_1}; // @[MSHR.scala 67:33]
  wire [7:0] _currentMask_T_1 = {io_from_addr_bits_tag_mask_7,io_from_addr_bits_tag_mask_6,io_from_addr_bits_tag_mask_5,
    io_from_addr_bits_tag_mask_4,io_from_addr_bits_tag_mask_3,io_from_addr_bits_tag_mask_2,io_from_addr_bits_tag_mask_1,
    io_from_addr_bits_tag_mask_0}; // @[MSHR.scala 70:70]
  wire [7:0] _GEN_56 = 2'h0 == valid_entry ? _currentMask_T_1 : currentMask_0; // @[MSHR.scala 24:28 70:{34,34}]
  wire [7:0] _GEN_57 = 2'h1 == valid_entry ? _currentMask_T_1 : currentMask_1; // @[MSHR.scala 24:28 70:{34,34}]
  wire [7:0] _GEN_58 = 2'h2 == valid_entry ? _currentMask_T_1 : currentMask_2; // @[MSHR.scala 24:28 70:{34,34}]
  wire [7:0] _GEN_59 = 2'h3 == valid_entry ? _currentMask_T_1 : currentMask_3; // @[MSHR.scala 24:28 70:{34,34}]
  wire  _GEN_127 = _T_1 ? 1'h0 : _io_idx_entry_T; // @[MSHR.scala 22:16 59:32]
  wire  _T_25 = 2'h1 == state; // @[MSHR.scala 57:16]
  wire [7:0] _currentMask_T_2 = {reg_req_mask_7,reg_req_mask_6,reg_req_mask_5,reg_req_mask_4,reg_req_mask_3,
    reg_req_mask_2,reg_req_mask_1,reg_req_mask_0}; // @[MSHR.scala 80:48]
  wire  _T_28 = io_to_pipe_ready & io_to_pipe_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _used_T_12 = 4'h1 << output_entry; // @[MSHR.scala 83:48]
  wire [3:0] _used_T_15 = _valid_entry_T_1 | _used_T_12; // @[MSHR.scala 83:48]
  wire [3:0] _used_T_16 = ~_used_T_15; // @[MSHR.scala 83:48]
  wire [3:0] _GEN_142 = _T_28 ? _used_T_16 : used; // @[MSHR.scala 26:21 83:{28,34}]
  wire [51:0] _output_tag_WIRE = tag_output_tag_MPORT_data;
  wire  output_tag_isWrite = _output_tag_WIRE[0]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_0 = _output_tag_WIRE[4:1]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_1 = _output_tag_WIRE[8:5]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_2 = _output_tag_WIRE[12:9]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_3 = _output_tag_WIRE[16:13]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_4 = _output_tag_WIRE[20:17]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_5 = _output_tag_WIRE[24:21]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_6 = _output_tag_WIRE[28:25]; // @[MSHR.scala 86:51]
  wire [3:0] output_tag_wordOffset1H_7 = _output_tag_WIRE[32:29]; // @[MSHR.scala 86:51]
  wire  output_tag_isvec = _output_tag_WIRE[33]; // @[MSHR.scala 86:51]
  wire  output_tag_unsigned = _output_tag_WIRE[34]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_0 = _output_tag_WIRE[35]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_1 = _output_tag_WIRE[36]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_2 = _output_tag_WIRE[37]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_3 = _output_tag_WIRE[38]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_4 = _output_tag_WIRE[39]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_5 = _output_tag_WIRE[40]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_6 = _output_tag_WIRE[41]; // @[MSHR.scala 86:51]
  wire  output_tag_mask_7 = _output_tag_WIRE[42]; // @[MSHR.scala 86:51]
  wire [4:0] output_tag_reg_idxw = _output_tag_WIRE[47:43]; // @[MSHR.scala 86:51]
  wire  output_tag_wxd = _output_tag_WIRE[48]; // @[MSHR.scala 86:51]
  wire  output_tag_wfd = _output_tag_WIRE[49]; // @[MSHR.scala 86:51]
  wire [1:0] output_tag_warp_id = _output_tag_WIRE[51:50]; // @[MSHR.scala 86:51]
  wire  _output_data_0_result_T = output_tag_wordOffset1H_0 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_0_result_T_1 = output_tag_wordOffset1H_0 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_0_result_T_4 = ~data_0_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_0_result_T_6 = {16'h0,data_0_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_8 = {16'hffff,data_0_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_9 = ~data_0_raw_data_data[31] | output_tag_unsigned ? _output_data_0_result_T_6 :
    _output_data_0_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_0_result_T_10 = output_tag_wordOffset1H_0 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_0_result_T_13 = ~data_0_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_0_result_T_15 = {16'h0,data_0_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_17 = {16'hffff,data_0_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_18 = ~data_0_raw_data_data[15] | output_tag_unsigned ? _output_data_0_result_T_15
     : _output_data_0_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_0_result_T_19 = output_tag_wordOffset1H_0 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_0_result_T_24 = {24'h0,data_0_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_26 = {24'hffffff,data_0_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_27 = _output_data_0_result_T_4 ? _output_data_0_result_T_24 :
    _output_data_0_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_0_result_T_28 = output_tag_wordOffset1H_0 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_0_result_T_33 = {24'h0,data_0_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_35 = {24'hffffff,data_0_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_36 = ~data_0_raw_data_data[23] | output_tag_unsigned ? _output_data_0_result_T_33
     : _output_data_0_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_0_result_T_37 = output_tag_wordOffset1H_0 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_0_result_T_42 = {24'h0,data_0_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_44 = {24'hffffff,data_0_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_45 = _output_data_0_result_T_13 ? _output_data_0_result_T_42 :
    _output_data_0_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_0_result_T_46 = output_tag_wordOffset1H_0 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_0_result_T_51 = {24'h0,data_0_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_53 = {24'hffffff,data_0_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_0_result_T_54 = ~data_0_raw_data_data[7] | output_tag_unsigned ? _output_data_0_result_T_51
     : _output_data_0_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_0_result_T_55 = _output_data_0_result_T_46 ? _output_data_0_result_T_54 :
    data_0_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_0_result_T_56 = _output_data_0_result_T_37 ? _output_data_0_result_T_45 :
    _output_data_0_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_0_result_T_57 = _output_data_0_result_T_28 ? _output_data_0_result_T_36 :
    _output_data_0_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_0_result_T_58 = _output_data_0_result_T_19 ? _output_data_0_result_T_27 :
    _output_data_0_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_0_result_T_59 = _output_data_0_result_T_10 ? _output_data_0_result_T_18 :
    _output_data_0_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_0_result_T_60 = _output_data_0_result_T_1 ? _output_data_0_result_T_9 :
    _output_data_0_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_0_result = _output_data_0_result_T ? data_0_raw_data_data : _output_data_0_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_1_result_T = output_tag_wordOffset1H_1 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_1_result_T_1 = output_tag_wordOffset1H_1 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_1_result_T_4 = ~data_1_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_1_result_T_6 = {16'h0,data_1_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_8 = {16'hffff,data_1_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_9 = ~data_1_raw_data_data[31] | output_tag_unsigned ? _output_data_1_result_T_6 :
    _output_data_1_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_1_result_T_10 = output_tag_wordOffset1H_1 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_1_result_T_13 = ~data_1_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_1_result_T_15 = {16'h0,data_1_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_17 = {16'hffff,data_1_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_18 = ~data_1_raw_data_data[15] | output_tag_unsigned ? _output_data_1_result_T_15
     : _output_data_1_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_1_result_T_19 = output_tag_wordOffset1H_1 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_1_result_T_24 = {24'h0,data_1_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_26 = {24'hffffff,data_1_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_27 = _output_data_1_result_T_4 ? _output_data_1_result_T_24 :
    _output_data_1_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_1_result_T_28 = output_tag_wordOffset1H_1 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_1_result_T_33 = {24'h0,data_1_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_35 = {24'hffffff,data_1_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_36 = ~data_1_raw_data_data[23] | output_tag_unsigned ? _output_data_1_result_T_33
     : _output_data_1_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_1_result_T_37 = output_tag_wordOffset1H_1 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_1_result_T_42 = {24'h0,data_1_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_44 = {24'hffffff,data_1_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_45 = _output_data_1_result_T_13 ? _output_data_1_result_T_42 :
    _output_data_1_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_1_result_T_46 = output_tag_wordOffset1H_1 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_1_result_T_51 = {24'h0,data_1_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_53 = {24'hffffff,data_1_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_1_result_T_54 = ~data_1_raw_data_data[7] | output_tag_unsigned ? _output_data_1_result_T_51
     : _output_data_1_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_1_result_T_55 = _output_data_1_result_T_46 ? _output_data_1_result_T_54 :
    data_1_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_1_result_T_56 = _output_data_1_result_T_37 ? _output_data_1_result_T_45 :
    _output_data_1_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_1_result_T_57 = _output_data_1_result_T_28 ? _output_data_1_result_T_36 :
    _output_data_1_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_1_result_T_58 = _output_data_1_result_T_19 ? _output_data_1_result_T_27 :
    _output_data_1_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_1_result_T_59 = _output_data_1_result_T_10 ? _output_data_1_result_T_18 :
    _output_data_1_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_1_result_T_60 = _output_data_1_result_T_1 ? _output_data_1_result_T_9 :
    _output_data_1_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_1_result = _output_data_1_result_T ? data_1_raw_data_data : _output_data_1_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_2_result_T = output_tag_wordOffset1H_2 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_2_result_T_1 = output_tag_wordOffset1H_2 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_2_result_T_4 = ~data_2_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_2_result_T_6 = {16'h0,data_2_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_8 = {16'hffff,data_2_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_9 = ~data_2_raw_data_data[31] | output_tag_unsigned ? _output_data_2_result_T_6 :
    _output_data_2_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_2_result_T_10 = output_tag_wordOffset1H_2 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_2_result_T_13 = ~data_2_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_2_result_T_15 = {16'h0,data_2_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_17 = {16'hffff,data_2_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_18 = ~data_2_raw_data_data[15] | output_tag_unsigned ? _output_data_2_result_T_15
     : _output_data_2_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_2_result_T_19 = output_tag_wordOffset1H_2 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_2_result_T_24 = {24'h0,data_2_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_26 = {24'hffffff,data_2_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_27 = _output_data_2_result_T_4 ? _output_data_2_result_T_24 :
    _output_data_2_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_2_result_T_28 = output_tag_wordOffset1H_2 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_2_result_T_33 = {24'h0,data_2_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_35 = {24'hffffff,data_2_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_36 = ~data_2_raw_data_data[23] | output_tag_unsigned ? _output_data_2_result_T_33
     : _output_data_2_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_2_result_T_37 = output_tag_wordOffset1H_2 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_2_result_T_42 = {24'h0,data_2_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_44 = {24'hffffff,data_2_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_45 = _output_data_2_result_T_13 ? _output_data_2_result_T_42 :
    _output_data_2_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_2_result_T_46 = output_tag_wordOffset1H_2 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_2_result_T_51 = {24'h0,data_2_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_53 = {24'hffffff,data_2_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_2_result_T_54 = ~data_2_raw_data_data[7] | output_tag_unsigned ? _output_data_2_result_T_51
     : _output_data_2_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_2_result_T_55 = _output_data_2_result_T_46 ? _output_data_2_result_T_54 :
    data_2_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_2_result_T_56 = _output_data_2_result_T_37 ? _output_data_2_result_T_45 :
    _output_data_2_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_2_result_T_57 = _output_data_2_result_T_28 ? _output_data_2_result_T_36 :
    _output_data_2_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_2_result_T_58 = _output_data_2_result_T_19 ? _output_data_2_result_T_27 :
    _output_data_2_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_2_result_T_59 = _output_data_2_result_T_10 ? _output_data_2_result_T_18 :
    _output_data_2_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_2_result_T_60 = _output_data_2_result_T_1 ? _output_data_2_result_T_9 :
    _output_data_2_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_2_result = _output_data_2_result_T ? data_2_raw_data_data : _output_data_2_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_3_result_T = output_tag_wordOffset1H_3 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_3_result_T_1 = output_tag_wordOffset1H_3 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_3_result_T_4 = ~data_3_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_3_result_T_6 = {16'h0,data_3_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_8 = {16'hffff,data_3_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_9 = ~data_3_raw_data_data[31] | output_tag_unsigned ? _output_data_3_result_T_6 :
    _output_data_3_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_3_result_T_10 = output_tag_wordOffset1H_3 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_3_result_T_13 = ~data_3_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_3_result_T_15 = {16'h0,data_3_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_17 = {16'hffff,data_3_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_18 = ~data_3_raw_data_data[15] | output_tag_unsigned ? _output_data_3_result_T_15
     : _output_data_3_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_3_result_T_19 = output_tag_wordOffset1H_3 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_3_result_T_24 = {24'h0,data_3_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_26 = {24'hffffff,data_3_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_27 = _output_data_3_result_T_4 ? _output_data_3_result_T_24 :
    _output_data_3_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_3_result_T_28 = output_tag_wordOffset1H_3 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_3_result_T_33 = {24'h0,data_3_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_35 = {24'hffffff,data_3_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_36 = ~data_3_raw_data_data[23] | output_tag_unsigned ? _output_data_3_result_T_33
     : _output_data_3_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_3_result_T_37 = output_tag_wordOffset1H_3 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_3_result_T_42 = {24'h0,data_3_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_44 = {24'hffffff,data_3_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_45 = _output_data_3_result_T_13 ? _output_data_3_result_T_42 :
    _output_data_3_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_3_result_T_46 = output_tag_wordOffset1H_3 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_3_result_T_51 = {24'h0,data_3_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_53 = {24'hffffff,data_3_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_3_result_T_54 = ~data_3_raw_data_data[7] | output_tag_unsigned ? _output_data_3_result_T_51
     : _output_data_3_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_3_result_T_55 = _output_data_3_result_T_46 ? _output_data_3_result_T_54 :
    data_3_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_3_result_T_56 = _output_data_3_result_T_37 ? _output_data_3_result_T_45 :
    _output_data_3_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_3_result_T_57 = _output_data_3_result_T_28 ? _output_data_3_result_T_36 :
    _output_data_3_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_3_result_T_58 = _output_data_3_result_T_19 ? _output_data_3_result_T_27 :
    _output_data_3_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_3_result_T_59 = _output_data_3_result_T_10 ? _output_data_3_result_T_18 :
    _output_data_3_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_3_result_T_60 = _output_data_3_result_T_1 ? _output_data_3_result_T_9 :
    _output_data_3_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_3_result = _output_data_3_result_T ? data_3_raw_data_data : _output_data_3_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_4_result_T = output_tag_wordOffset1H_4 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_4_result_T_1 = output_tag_wordOffset1H_4 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_4_result_T_4 = ~data_4_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_4_result_T_6 = {16'h0,data_4_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_8 = {16'hffff,data_4_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_9 = ~data_4_raw_data_data[31] | output_tag_unsigned ? _output_data_4_result_T_6 :
    _output_data_4_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_4_result_T_10 = output_tag_wordOffset1H_4 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_4_result_T_13 = ~data_4_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_4_result_T_15 = {16'h0,data_4_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_17 = {16'hffff,data_4_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_18 = ~data_4_raw_data_data[15] | output_tag_unsigned ? _output_data_4_result_T_15
     : _output_data_4_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_4_result_T_19 = output_tag_wordOffset1H_4 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_4_result_T_24 = {24'h0,data_4_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_26 = {24'hffffff,data_4_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_27 = _output_data_4_result_T_4 ? _output_data_4_result_T_24 :
    _output_data_4_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_4_result_T_28 = output_tag_wordOffset1H_4 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_4_result_T_33 = {24'h0,data_4_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_35 = {24'hffffff,data_4_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_36 = ~data_4_raw_data_data[23] | output_tag_unsigned ? _output_data_4_result_T_33
     : _output_data_4_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_4_result_T_37 = output_tag_wordOffset1H_4 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_4_result_T_42 = {24'h0,data_4_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_44 = {24'hffffff,data_4_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_45 = _output_data_4_result_T_13 ? _output_data_4_result_T_42 :
    _output_data_4_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_4_result_T_46 = output_tag_wordOffset1H_4 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_4_result_T_51 = {24'h0,data_4_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_53 = {24'hffffff,data_4_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_4_result_T_54 = ~data_4_raw_data_data[7] | output_tag_unsigned ? _output_data_4_result_T_51
     : _output_data_4_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_4_result_T_55 = _output_data_4_result_T_46 ? _output_data_4_result_T_54 :
    data_4_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_4_result_T_56 = _output_data_4_result_T_37 ? _output_data_4_result_T_45 :
    _output_data_4_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_4_result_T_57 = _output_data_4_result_T_28 ? _output_data_4_result_T_36 :
    _output_data_4_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_4_result_T_58 = _output_data_4_result_T_19 ? _output_data_4_result_T_27 :
    _output_data_4_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_4_result_T_59 = _output_data_4_result_T_10 ? _output_data_4_result_T_18 :
    _output_data_4_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_4_result_T_60 = _output_data_4_result_T_1 ? _output_data_4_result_T_9 :
    _output_data_4_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_4_result = _output_data_4_result_T ? data_4_raw_data_data : _output_data_4_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_5_result_T = output_tag_wordOffset1H_5 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_5_result_T_1 = output_tag_wordOffset1H_5 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_5_result_T_4 = ~data_5_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_5_result_T_6 = {16'h0,data_5_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_8 = {16'hffff,data_5_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_9 = ~data_5_raw_data_data[31] | output_tag_unsigned ? _output_data_5_result_T_6 :
    _output_data_5_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_5_result_T_10 = output_tag_wordOffset1H_5 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_5_result_T_13 = ~data_5_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_5_result_T_15 = {16'h0,data_5_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_17 = {16'hffff,data_5_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_18 = ~data_5_raw_data_data[15] | output_tag_unsigned ? _output_data_5_result_T_15
     : _output_data_5_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_5_result_T_19 = output_tag_wordOffset1H_5 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_5_result_T_24 = {24'h0,data_5_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_26 = {24'hffffff,data_5_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_27 = _output_data_5_result_T_4 ? _output_data_5_result_T_24 :
    _output_data_5_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_5_result_T_28 = output_tag_wordOffset1H_5 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_5_result_T_33 = {24'h0,data_5_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_35 = {24'hffffff,data_5_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_36 = ~data_5_raw_data_data[23] | output_tag_unsigned ? _output_data_5_result_T_33
     : _output_data_5_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_5_result_T_37 = output_tag_wordOffset1H_5 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_5_result_T_42 = {24'h0,data_5_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_44 = {24'hffffff,data_5_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_45 = _output_data_5_result_T_13 ? _output_data_5_result_T_42 :
    _output_data_5_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_5_result_T_46 = output_tag_wordOffset1H_5 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_5_result_T_51 = {24'h0,data_5_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_53 = {24'hffffff,data_5_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_5_result_T_54 = ~data_5_raw_data_data[7] | output_tag_unsigned ? _output_data_5_result_T_51
     : _output_data_5_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_5_result_T_55 = _output_data_5_result_T_46 ? _output_data_5_result_T_54 :
    data_5_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_5_result_T_56 = _output_data_5_result_T_37 ? _output_data_5_result_T_45 :
    _output_data_5_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_5_result_T_57 = _output_data_5_result_T_28 ? _output_data_5_result_T_36 :
    _output_data_5_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_5_result_T_58 = _output_data_5_result_T_19 ? _output_data_5_result_T_27 :
    _output_data_5_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_5_result_T_59 = _output_data_5_result_T_10 ? _output_data_5_result_T_18 :
    _output_data_5_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_5_result_T_60 = _output_data_5_result_T_1 ? _output_data_5_result_T_9 :
    _output_data_5_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_5_result = _output_data_5_result_T ? data_5_raw_data_data : _output_data_5_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_6_result_T = output_tag_wordOffset1H_6 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_6_result_T_1 = output_tag_wordOffset1H_6 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_6_result_T_4 = ~data_6_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_6_result_T_6 = {16'h0,data_6_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_8 = {16'hffff,data_6_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_9 = ~data_6_raw_data_data[31] | output_tag_unsigned ? _output_data_6_result_T_6 :
    _output_data_6_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_6_result_T_10 = output_tag_wordOffset1H_6 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_6_result_T_13 = ~data_6_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_6_result_T_15 = {16'h0,data_6_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_17 = {16'hffff,data_6_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_18 = ~data_6_raw_data_data[15] | output_tag_unsigned ? _output_data_6_result_T_15
     : _output_data_6_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_6_result_T_19 = output_tag_wordOffset1H_6 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_6_result_T_24 = {24'h0,data_6_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_26 = {24'hffffff,data_6_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_27 = _output_data_6_result_T_4 ? _output_data_6_result_T_24 :
    _output_data_6_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_6_result_T_28 = output_tag_wordOffset1H_6 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_6_result_T_33 = {24'h0,data_6_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_35 = {24'hffffff,data_6_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_36 = ~data_6_raw_data_data[23] | output_tag_unsigned ? _output_data_6_result_T_33
     : _output_data_6_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_6_result_T_37 = output_tag_wordOffset1H_6 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_6_result_T_42 = {24'h0,data_6_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_44 = {24'hffffff,data_6_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_45 = _output_data_6_result_T_13 ? _output_data_6_result_T_42 :
    _output_data_6_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_6_result_T_46 = output_tag_wordOffset1H_6 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_6_result_T_51 = {24'h0,data_6_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_53 = {24'hffffff,data_6_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_6_result_T_54 = ~data_6_raw_data_data[7] | output_tag_unsigned ? _output_data_6_result_T_51
     : _output_data_6_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_6_result_T_55 = _output_data_6_result_T_46 ? _output_data_6_result_T_54 :
    data_6_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_6_result_T_56 = _output_data_6_result_T_37 ? _output_data_6_result_T_45 :
    _output_data_6_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_6_result_T_57 = _output_data_6_result_T_28 ? _output_data_6_result_T_36 :
    _output_data_6_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_6_result_T_58 = _output_data_6_result_T_19 ? _output_data_6_result_T_27 :
    _output_data_6_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_6_result_T_59 = _output_data_6_result_T_10 ? _output_data_6_result_T_18 :
    _output_data_6_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_6_result_T_60 = _output_data_6_result_T_1 ? _output_data_6_result_T_9 :
    _output_data_6_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_6_result = _output_data_6_result_T ? data_6_raw_data_data : _output_data_6_result_T_60; // @[Mux.scala 101:16]
  wire  _output_data_7_result_T = output_tag_wordOffset1H_7 == 4'hf; // @[LSU.scala 106:13]
  wire  _output_data_7_result_T_1 = output_tag_wordOffset1H_7 == 4'hc; // @[LSU.scala 107:13]
  wire  _output_data_7_result_T_4 = ~data_7_raw_data_data[31] | output_tag_unsigned; // @[LSU.scala 107:38]
  wire [31:0] _output_data_7_result_T_6 = {16'h0,data_7_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_8 = {16'hffff,data_7_raw_data_data[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_9 = ~data_7_raw_data_data[31] | output_tag_unsigned ? _output_data_7_result_T_6 :
    _output_data_7_result_T_8; // @[LSU.scala 107:30]
  wire  _output_data_7_result_T_10 = output_tag_wordOffset1H_7 == 4'h3; // @[LSU.scala 108:13]
  wire  _output_data_7_result_T_13 = ~data_7_raw_data_data[15] | output_tag_unsigned; // @[LSU.scala 108:38]
  wire [31:0] _output_data_7_result_T_15 = {16'h0,data_7_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_17 = {16'hffff,data_7_raw_data_data[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_18 = ~data_7_raw_data_data[15] | output_tag_unsigned ? _output_data_7_result_T_15
     : _output_data_7_result_T_17; // @[LSU.scala 108:30]
  wire  _output_data_7_result_T_19 = output_tag_wordOffset1H_7 == 4'h8; // @[LSU.scala 109:13]
  wire [31:0] _output_data_7_result_T_24 = {24'h0,data_7_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_26 = {24'hffffff,data_7_raw_data_data[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_27 = _output_data_7_result_T_4 ? _output_data_7_result_T_24 :
    _output_data_7_result_T_26; // @[LSU.scala 109:30]
  wire  _output_data_7_result_T_28 = output_tag_wordOffset1H_7 == 4'h4; // @[LSU.scala 110:13]
  wire [31:0] _output_data_7_result_T_33 = {24'h0,data_7_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_35 = {24'hffffff,data_7_raw_data_data[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_36 = ~data_7_raw_data_data[23] | output_tag_unsigned ? _output_data_7_result_T_33
     : _output_data_7_result_T_35; // @[LSU.scala 110:30]
  wire  _output_data_7_result_T_37 = output_tag_wordOffset1H_7 == 4'h2; // @[LSU.scala 111:13]
  wire [31:0] _output_data_7_result_T_42 = {24'h0,data_7_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_44 = {24'hffffff,data_7_raw_data_data[15:8]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_45 = _output_data_7_result_T_13 ? _output_data_7_result_T_42 :
    _output_data_7_result_T_44; // @[LSU.scala 111:30]
  wire  _output_data_7_result_T_46 = output_tag_wordOffset1H_7 == 4'h1; // @[LSU.scala 112:13]
  wire [31:0] _output_data_7_result_T_51 = {24'h0,data_7_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_53 = {24'hffffff,data_7_raw_data_data[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _output_data_7_result_T_54 = ~data_7_raw_data_data[7] | output_tag_unsigned ? _output_data_7_result_T_51
     : _output_data_7_result_T_53; // @[LSU.scala 112:30]
  wire [31:0] _output_data_7_result_T_55 = _output_data_7_result_T_46 ? _output_data_7_result_T_54 :
    data_7_raw_data_data; // @[Mux.scala 101:16]
  wire [31:0] _output_data_7_result_T_56 = _output_data_7_result_T_37 ? _output_data_7_result_T_45 :
    _output_data_7_result_T_55; // @[Mux.scala 101:16]
  wire [31:0] _output_data_7_result_T_57 = _output_data_7_result_T_28 ? _output_data_7_result_T_36 :
    _output_data_7_result_T_56; // @[Mux.scala 101:16]
  wire [31:0] _output_data_7_result_T_58 = _output_data_7_result_T_19 ? _output_data_7_result_T_27 :
    _output_data_7_result_T_57; // @[Mux.scala 101:16]
  wire [31:0] _output_data_7_result_T_59 = _output_data_7_result_T_10 ? _output_data_7_result_T_18 :
    _output_data_7_result_T_58; // @[Mux.scala 101:16]
  wire [31:0] _output_data_7_result_T_60 = _output_data_7_result_T_1 ? _output_data_7_result_T_9 :
    _output_data_7_result_T_59; // @[Mux.scala 101:16]
  wire [31:0] output_data_7_result = _output_data_7_result_T ? data_7_raw_data_data : _output_data_7_result_T_60; // @[Mux.scala 101:16]
  wire [16:0] io_to_pipe_bits_tag_lo_lo = {output_tag_wordOffset1H_3,output_tag_wordOffset1H_2,output_tag_wordOffset1H_1
    ,output_tag_wordOffset1H_0,output_tag_isWrite}; // @[MSHR.scala 96:45]
  wire [34:0] io_to_pipe_bits_tag_lo = {output_tag_unsigned,output_tag_isvec,output_tag_wordOffset1H_7,
    output_tag_wordOffset1H_6,output_tag_wordOffset1H_5,output_tag_wordOffset1H_4,io_to_pipe_bits_tag_lo_lo}; // @[MSHR.scala 96:45]
  wire [5:0] io_to_pipe_bits_tag_hi_lo = {output_tag_mask_5,output_tag_mask_4,output_tag_mask_3,output_tag_mask_2,
    output_tag_mask_1,output_tag_mask_0}; // @[MSHR.scala 96:45]
  wire [51:0] _io_to_pipe_bits_tag_T = {output_tag_warp_id,output_tag_wfd,output_tag_wxd,output_tag_reg_idxw,
    output_tag_mask_7,output_tag_mask_6,io_to_pipe_bits_tag_hi_lo,io_to_pipe_bits_tag_lo}; // @[MSHR.scala 96:45]
  assign data_0_raw_data_en = 1'h1;
  assign data_0_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_0_raw_data_data = data_0[data_0_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_0_MPORT_data = io_from_dcache_bits_data_0;
  assign data_0_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_0_MPORT_mask = io_from_dcache_bits_activeMask_0;
  assign data_0_MPORT_en = _T_20 & _T_1;
  assign data_0_MPORT_2_data = 32'h0;
  assign data_0_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_0_MPORT_2_mask = 1'h1;
  assign data_0_MPORT_2_en = _T_20 & _GEN_127;
  assign data_0_MPORT_4_data = 32'h0;
  assign data_0_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_0_MPORT_4_mask = 1'h1;
  assign data_0_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_1_raw_data_en = 1'h1;
  assign data_1_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_1_raw_data_data = data_1[data_1_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_1_MPORT_data = io_from_dcache_bits_data_1;
  assign data_1_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_1_MPORT_mask = io_from_dcache_bits_activeMask_1;
  assign data_1_MPORT_en = _T_20 & _T_1;
  assign data_1_MPORT_2_data = 32'h0;
  assign data_1_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_1_MPORT_2_mask = 1'h1;
  assign data_1_MPORT_2_en = _T_20 & _GEN_127;
  assign data_1_MPORT_4_data = 32'h0;
  assign data_1_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_1_MPORT_4_mask = 1'h1;
  assign data_1_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_2_raw_data_en = 1'h1;
  assign data_2_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_2_raw_data_data = data_2[data_2_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_2_MPORT_data = io_from_dcache_bits_data_2;
  assign data_2_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_2_MPORT_mask = io_from_dcache_bits_activeMask_2;
  assign data_2_MPORT_en = _T_20 & _T_1;
  assign data_2_MPORT_2_data = 32'h0;
  assign data_2_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_2_MPORT_2_mask = 1'h1;
  assign data_2_MPORT_2_en = _T_20 & _GEN_127;
  assign data_2_MPORT_4_data = 32'h0;
  assign data_2_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_2_MPORT_4_mask = 1'h1;
  assign data_2_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_3_raw_data_en = 1'h1;
  assign data_3_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_3_raw_data_data = data_3[data_3_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_3_MPORT_data = io_from_dcache_bits_data_3;
  assign data_3_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_3_MPORT_mask = io_from_dcache_bits_activeMask_3;
  assign data_3_MPORT_en = _T_20 & _T_1;
  assign data_3_MPORT_2_data = 32'h0;
  assign data_3_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_3_MPORT_2_mask = 1'h1;
  assign data_3_MPORT_2_en = _T_20 & _GEN_127;
  assign data_3_MPORT_4_data = 32'h0;
  assign data_3_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_3_MPORT_4_mask = 1'h1;
  assign data_3_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_4_raw_data_en = 1'h1;
  assign data_4_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_4_raw_data_data = data_4[data_4_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_4_MPORT_data = io_from_dcache_bits_data_4;
  assign data_4_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_4_MPORT_mask = io_from_dcache_bits_activeMask_4;
  assign data_4_MPORT_en = _T_20 & _T_1;
  assign data_4_MPORT_2_data = 32'h0;
  assign data_4_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_4_MPORT_2_mask = 1'h1;
  assign data_4_MPORT_2_en = _T_20 & _GEN_127;
  assign data_4_MPORT_4_data = 32'h0;
  assign data_4_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_4_MPORT_4_mask = 1'h1;
  assign data_4_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_5_raw_data_en = 1'h1;
  assign data_5_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_5_raw_data_data = data_5[data_5_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_5_MPORT_data = io_from_dcache_bits_data_5;
  assign data_5_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_5_MPORT_mask = io_from_dcache_bits_activeMask_5;
  assign data_5_MPORT_en = _T_20 & _T_1;
  assign data_5_MPORT_2_data = 32'h0;
  assign data_5_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_5_MPORT_2_mask = 1'h1;
  assign data_5_MPORT_2_en = _T_20 & _GEN_127;
  assign data_5_MPORT_4_data = 32'h0;
  assign data_5_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_5_MPORT_4_mask = 1'h1;
  assign data_5_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_6_raw_data_en = 1'h1;
  assign data_6_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_6_raw_data_data = data_6[data_6_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_6_MPORT_data = io_from_dcache_bits_data_6;
  assign data_6_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_6_MPORT_mask = io_from_dcache_bits_activeMask_6;
  assign data_6_MPORT_en = _T_20 & _T_1;
  assign data_6_MPORT_2_data = 32'h0;
  assign data_6_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_6_MPORT_2_mask = 1'h1;
  assign data_6_MPORT_2_en = _T_20 & _GEN_127;
  assign data_6_MPORT_4_data = 32'h0;
  assign data_6_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_6_MPORT_4_mask = 1'h1;
  assign data_6_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign data_7_raw_data_en = 1'h1;
  assign data_7_raw_data_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign data_7_raw_data_data = data_7[data_7_raw_data_addr]; // @[MSHR.scala 21:17]
  assign data_7_MPORT_data = io_from_dcache_bits_data_7;
  assign data_7_MPORT_addr = io_from_dcache_bits_instrId;
  assign data_7_MPORT_mask = io_from_dcache_bits_activeMask_7;
  assign data_7_MPORT_en = _T_20 & _T_1;
  assign data_7_MPORT_2_data = 32'h0;
  assign data_7_MPORT_2_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_7_MPORT_2_mask = 1'h1;
  assign data_7_MPORT_2_en = _T_20 & _GEN_127;
  assign data_7_MPORT_4_data = 32'h0;
  assign data_7_MPORT_4_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign data_7_MPORT_4_mask = 1'h1;
  assign data_7_MPORT_4_en = _T_20 ? 1'h0 : _T_25;
  assign tag_output_tag_MPORT_en = 1'h1;
  assign tag_output_tag_MPORT_addr = _output_entry_T ? _output_entry_T_7 : 2'h0;
  assign tag_output_tag_MPORT_data = tag[tag_output_tag_MPORT_addr]; // @[MSHR.scala 22:16]
  assign tag_MPORT_1_data = {hi_1,lo_1};
  assign tag_MPORT_1_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign tag_MPORT_1_mask = 1'h1;
  assign tag_MPORT_1_en = _T_20 & _GEN_127;
  assign tag_MPORT_3_data = {hi_1,lo_1};
  assign tag_MPORT_3_addr = _valid_entry_T ? 2'h0 : _valid_entry_T_8;
  assign tag_MPORT_3_mask = 1'h1;
  assign tag_MPORT_3_en = _T_20 ? 1'h0 : _T_25;
  assign io_from_addr_ready = _io_from_dcache_ready_T & ~_valid_entry_T; // @[MSHR.scala 36:40]
  assign io_idx_entry = _io_idx_entry_T ? valid_entry : 2'h0; // @[MSHR.scala 37:22]
  assign io_from_dcache_ready = state == 2'h0; // @[MSHR.scala 35:32]
  assign io_to_pipe_valid = _output_entry_T & _T_8; // @[MSHR.scala 95:36]
  assign io_to_pipe_bits_tag_warp_id = _io_to_pipe_bits_tag_T[51:50]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_wfd = _io_to_pipe_bits_tag_T[49]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_wxd = _io_to_pipe_bits_tag_T[48]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_reg_idxw = _io_to_pipe_bits_tag_T[47:43]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_0 = _io_to_pipe_bits_tag_T[35]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_1 = _io_to_pipe_bits_tag_T[36]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_2 = _io_to_pipe_bits_tag_T[37]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_3 = _io_to_pipe_bits_tag_T[38]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_4 = _io_to_pipe_bits_tag_T[39]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_5 = _io_to_pipe_bits_tag_T[40]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_6 = _io_to_pipe_bits_tag_T[41]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_mask_7 = _io_to_pipe_bits_tag_T[42]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_tag_isWrite = _io_to_pipe_bits_tag_T[0]; // @[MSHR.scala 96:45]
  assign io_to_pipe_bits_data_0 = output_tag_mask_0 ? output_data_0_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_1 = output_tag_mask_1 ? output_data_1_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_2 = output_tag_mask_2 ? output_data_2_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_3 = output_tag_mask_3 ? output_data_3_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_4 = output_tag_mask_4 ? output_data_4_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_5 = output_tag_mask_5 ? output_data_5_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_6 = output_tag_mask_6 ? output_data_6_result : 32'h0; // @[MSHR.scala 90:26]
  assign io_to_pipe_bits_data_7 = output_tag_mask_7 ? output_data_7_result : 32'h0; // @[MSHR.scala 90:26]
  always @(posedge clock) begin
    if (data_0_MPORT_en & data_0_MPORT_mask) begin
      data_0[data_0_MPORT_addr] <= data_0_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_0_MPORT_2_en & data_0_MPORT_2_mask) begin
      data_0[data_0_MPORT_2_addr] <= data_0_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_0_MPORT_4_en & data_0_MPORT_4_mask) begin
      data_0[data_0_MPORT_4_addr] <= data_0_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_1_MPORT_en & data_1_MPORT_mask) begin
      data_1[data_1_MPORT_addr] <= data_1_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_1_MPORT_2_en & data_1_MPORT_2_mask) begin
      data_1[data_1_MPORT_2_addr] <= data_1_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_1_MPORT_4_en & data_1_MPORT_4_mask) begin
      data_1[data_1_MPORT_4_addr] <= data_1_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_2_MPORT_en & data_2_MPORT_mask) begin
      data_2[data_2_MPORT_addr] <= data_2_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_2_MPORT_2_en & data_2_MPORT_2_mask) begin
      data_2[data_2_MPORT_2_addr] <= data_2_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_2_MPORT_4_en & data_2_MPORT_4_mask) begin
      data_2[data_2_MPORT_4_addr] <= data_2_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_3_MPORT_en & data_3_MPORT_mask) begin
      data_3[data_3_MPORT_addr] <= data_3_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_3_MPORT_2_en & data_3_MPORT_2_mask) begin
      data_3[data_3_MPORT_2_addr] <= data_3_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_3_MPORT_4_en & data_3_MPORT_4_mask) begin
      data_3[data_3_MPORT_4_addr] <= data_3_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_4_MPORT_en & data_4_MPORT_mask) begin
      data_4[data_4_MPORT_addr] <= data_4_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_4_MPORT_2_en & data_4_MPORT_2_mask) begin
      data_4[data_4_MPORT_2_addr] <= data_4_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_4_MPORT_4_en & data_4_MPORT_4_mask) begin
      data_4[data_4_MPORT_4_addr] <= data_4_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_5_MPORT_en & data_5_MPORT_mask) begin
      data_5[data_5_MPORT_addr] <= data_5_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_5_MPORT_2_en & data_5_MPORT_2_mask) begin
      data_5[data_5_MPORT_2_addr] <= data_5_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_5_MPORT_4_en & data_5_MPORT_4_mask) begin
      data_5[data_5_MPORT_4_addr] <= data_5_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_6_MPORT_en & data_6_MPORT_mask) begin
      data_6[data_6_MPORT_addr] <= data_6_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_6_MPORT_2_en & data_6_MPORT_2_mask) begin
      data_6[data_6_MPORT_2_addr] <= data_6_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_6_MPORT_4_en & data_6_MPORT_4_mask) begin
      data_6[data_6_MPORT_4_addr] <= data_6_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (data_7_MPORT_en & data_7_MPORT_mask) begin
      data_7[data_7_MPORT_addr] <= data_7_MPORT_data; // @[MSHR.scala 21:17]
    end
    if (data_7_MPORT_2_en & data_7_MPORT_2_mask) begin
      data_7[data_7_MPORT_2_addr] <= data_7_MPORT_2_data; // @[MSHR.scala 21:17]
    end
    if (data_7_MPORT_4_en & data_7_MPORT_4_mask) begin
      data_7[data_7_MPORT_4_addr] <= data_7_MPORT_4_data; // @[MSHR.scala 21:17]
    end
    if (tag_MPORT_1_en & tag_MPORT_1_mask) begin
      tag[tag_MPORT_1_addr] <= tag_MPORT_1_data; // @[MSHR.scala 22:16]
    end
    if (tag_MPORT_3_en & tag_MPORT_3_mask) begin
      tag[tag_MPORT_3_addr] <= tag_MPORT_3_data; // @[MSHR.scala 22:16]
    end
    if (reset) begin // @[MSHR.scala 24:28]
      currentMask_0 <= 8'h0; // @[MSHR.scala 24:28]
    end else if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (2'h0 == io_from_dcache_bits_instrId) begin // @[MSHR.scala 61:50]
          currentMask_0 <= _currentMask_T; // @[MSHR.scala 61:50]
        end
      end else if (_io_idx_entry_T) begin // @[MSHR.scala 63:36]
        currentMask_0 <= _GEN_56;
      end
    end else if (2'h1 == state) begin // @[MSHR.scala 57:16]
      if (2'h0 == valid_entry) begin // @[MSHR.scala 80:32]
        currentMask_0 <= _currentMask_T_2; // @[MSHR.scala 80:32]
      end
    end
    if (reset) begin // @[MSHR.scala 24:28]
      currentMask_1 <= 8'h0; // @[MSHR.scala 24:28]
    end else if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (2'h1 == io_from_dcache_bits_instrId) begin // @[MSHR.scala 61:50]
          currentMask_1 <= _currentMask_T; // @[MSHR.scala 61:50]
        end
      end else if (_io_idx_entry_T) begin // @[MSHR.scala 63:36]
        currentMask_1 <= _GEN_57;
      end
    end else if (2'h1 == state) begin // @[MSHR.scala 57:16]
      if (2'h1 == valid_entry) begin // @[MSHR.scala 80:32]
        currentMask_1 <= _currentMask_T_2; // @[MSHR.scala 80:32]
      end
    end
    if (reset) begin // @[MSHR.scala 24:28]
      currentMask_2 <= 8'h0; // @[MSHR.scala 24:28]
    end else if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (2'h2 == io_from_dcache_bits_instrId) begin // @[MSHR.scala 61:50]
          currentMask_2 <= _currentMask_T; // @[MSHR.scala 61:50]
        end
      end else if (_io_idx_entry_T) begin // @[MSHR.scala 63:36]
        currentMask_2 <= _GEN_58;
      end
    end else if (2'h1 == state) begin // @[MSHR.scala 57:16]
      if (2'h2 == valid_entry) begin // @[MSHR.scala 80:32]
        currentMask_2 <= _currentMask_T_2; // @[MSHR.scala 80:32]
      end
    end
    if (reset) begin // @[MSHR.scala 24:28]
      currentMask_3 <= 8'h0; // @[MSHR.scala 24:28]
    end else if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (2'h3 == io_from_dcache_bits_instrId) begin // @[MSHR.scala 61:50]
          currentMask_3 <= _currentMask_T; // @[MSHR.scala 61:50]
        end
      end else if (_io_idx_entry_T) begin // @[MSHR.scala 63:36]
        currentMask_3 <= _GEN_59;
      end
    end else if (2'h1 == state) begin // @[MSHR.scala 57:16]
      if (2'h3 == valid_entry) begin // @[MSHR.scala 80:32]
        currentMask_3 <= _currentMask_T_2; // @[MSHR.scala 80:32]
      end
    end
    if (reset) begin // @[MSHR.scala 26:21]
      used <= 4'h0; // @[MSHR.scala 26:21]
    end else if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (!(_T_1)) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 63:36]
          used <= _used_T_1; // @[MSHR.scala 64:14]
        end
      end
    end else if (2'h1 == state) begin // @[MSHR.scala 57:16]
      used <= _used_T_1; // @[MSHR.scala 74:12]
    end else if (2'h2 == state) begin // @[MSHR.scala 57:16]
      used <= _GEN_142;
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_0 <= io_from_addr_bits_tag_mask_0; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_1 <= io_from_addr_bits_tag_mask_1; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_2 <= io_from_addr_bits_tag_mask_2; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_3 <= io_from_addr_bits_tag_mask_3; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_4 <= io_from_addr_bits_tag_mask_4; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_5 <= io_from_addr_bits_tag_mask_5; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_6 <= io_from_addr_bits_tag_mask_6; // @[MSHR.scala 62:41]
        end
      end
    end
    if (2'h0 == state) begin // @[MSHR.scala 57:16]
      if (_T_1) begin // @[MSHR.scala 59:32]
        if (_io_idx_entry_T) begin // @[MSHR.scala 62:32]
          reg_req_mask_7 <= io_from_addr_bits_tag_mask_7; // @[MSHR.scala 62:41]
        end
      end
    end
    if (reset) begin // @[MSHR.scala 33:22]
      state <= 2'h0; // @[MSHR.scala 33:22]
    end else if (_io_from_dcache_ready_T) begin // @[MSHR.scala 39:23]
      if (_T_1) begin // @[MSHR.scala 40:30]
        if (_io_idx_entry_T) begin // @[MSHR.scala 41:30]
          state <= 2'h1; // @[MSHR.scala 42:15]
        end else begin
          state <= _GEN_4;
        end
      end else if (_output_entry_T & io_to_pipe_ready) begin // @[MSHR.scala 46:47]
        state <= 2'h2; // @[MSHR.scala 47:13]
      end else begin
        state <= 2'h0; // @[MSHR.scala 49:13]
      end
    end else if (state == 2'h2) begin // @[MSHR.scala 51:28]
      if (io_to_pipe_ready & |_T_13) begin // @[MSHR.scala 52:72]
        state <= 2'h2; // @[MSHR.scala 52:78]
      end else begin
        state <= 2'h0; // @[MSHR.scala 52:102]
      end
    end else if (state == 2'h1) begin // @[MSHR.scala 53:28]
      state <= _GEN_9;
    end else begin
      state <= 2'h0; // @[MSHR.scala 55:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_0[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_1[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_2[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_3[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_4[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_5[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_6[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data_7[initvar] = _RAND_7[31:0];
  _RAND_8 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    tag[initvar] = _RAND_8[51:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  currentMask_0 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  currentMask_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  currentMask_2 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  currentMask_3 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  used = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  reg_req_mask_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_req_mask_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  reg_req_mask_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reg_req_mask_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reg_req_mask_4 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  reg_req_mask_5 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  reg_req_mask_6 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  reg_req_mask_7 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  state = _RAND_22[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ShiftBoard(
  input   clock,
  input   reset,
  input   io_left,
  input   io_right,
  output  io_full,
  output  io_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  taps_0; // @[LSU.scala 373:36]
  reg  taps_1; // @[LSU.scala 373:36]
  reg  taps_2; // @[LSU.scala 373:36]
  reg  taps_3; // @[LSU.scala 373:36]
  wire  _taps_0_T = io_left ^ io_right; // @[LSU.scala 378:31]
  wire  _taps_0_T_2 = io_left ^ io_right ? io_left | taps_1 : taps_0; // @[LSU.scala 378:21]
  assign io_full = taps_3; // @[LSU.scala 382:10]
  assign io_empty = ~_taps_0_T_2; // @[LSU.scala 383:14]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 373:36]
      taps_0 <= 1'h0; // @[LSU.scala 373:36]
    end else if (io_left ^ io_right) begin // @[LSU.scala 378:21]
      taps_0 <= io_left | taps_1;
    end
    if (reset) begin // @[LSU.scala 373:36]
      taps_1 <= 1'h0; // @[LSU.scala 373:36]
    end else if (_taps_0_T) begin // @[LSU.scala 380:16]
      if (io_left) begin // @[LSU.scala 380:41]
        taps_1 <= taps_0;
      end else begin
        taps_1 <= taps_2;
      end
    end
    if (reset) begin // @[LSU.scala 373:36]
      taps_2 <= 1'h0; // @[LSU.scala 373:36]
    end else if (_taps_0_T) begin // @[LSU.scala 380:16]
      if (io_left) begin // @[LSU.scala 380:41]
        taps_2 <= taps_1;
      end else begin
        taps_2 <= taps_3;
      end
    end
    if (reset) begin // @[LSU.scala 373:36]
      taps_3 <= 1'h0; // @[LSU.scala 373:36]
    end else if (_taps_0_T) begin // @[LSU.scala 379:32]
      taps_3 <= io_left & taps_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  taps_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  taps_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  taps_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  taps_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSUexe(
  input         clock,
  input         reset,
  output        io_lsu_req_ready,
  input         io_lsu_req_valid,
  input  [31:0] io_lsu_req_bits_in1_0,
  input  [31:0] io_lsu_req_bits_in1_1,
  input  [31:0] io_lsu_req_bits_in1_2,
  input  [31:0] io_lsu_req_bits_in1_3,
  input  [31:0] io_lsu_req_bits_in1_4,
  input  [31:0] io_lsu_req_bits_in1_5,
  input  [31:0] io_lsu_req_bits_in1_6,
  input  [31:0] io_lsu_req_bits_in1_7,
  input  [31:0] io_lsu_req_bits_in2_0,
  input  [31:0] io_lsu_req_bits_in2_1,
  input  [31:0] io_lsu_req_bits_in2_2,
  input  [31:0] io_lsu_req_bits_in2_3,
  input  [31:0] io_lsu_req_bits_in2_4,
  input  [31:0] io_lsu_req_bits_in2_5,
  input  [31:0] io_lsu_req_bits_in2_6,
  input  [31:0] io_lsu_req_bits_in2_7,
  input  [31:0] io_lsu_req_bits_in3_0,
  input  [31:0] io_lsu_req_bits_in3_1,
  input  [31:0] io_lsu_req_bits_in3_2,
  input  [31:0] io_lsu_req_bits_in3_3,
  input  [31:0] io_lsu_req_bits_in3_4,
  input  [31:0] io_lsu_req_bits_in3_5,
  input  [31:0] io_lsu_req_bits_in3_6,
  input  [31:0] io_lsu_req_bits_in3_7,
  input         io_lsu_req_bits_mask_0,
  input         io_lsu_req_bits_mask_1,
  input         io_lsu_req_bits_mask_2,
  input         io_lsu_req_bits_mask_3,
  input         io_lsu_req_bits_mask_4,
  input         io_lsu_req_bits_mask_5,
  input         io_lsu_req_bits_mask_6,
  input         io_lsu_req_bits_mask_7,
  input  [31:0] io_lsu_req_bits_ctrl_inst,
  input  [1:0]  io_lsu_req_bits_ctrl_wid,
  input         io_lsu_req_bits_ctrl_fp,
  input  [1:0]  io_lsu_req_bits_ctrl_branch,
  input         io_lsu_req_bits_ctrl_simt_stack,
  input         io_lsu_req_bits_ctrl_simt_stack_op,
  input         io_lsu_req_bits_ctrl_barrier,
  input  [1:0]  io_lsu_req_bits_ctrl_csr,
  input         io_lsu_req_bits_ctrl_reverse,
  input         io_lsu_req_bits_ctrl_isvec,
  input         io_lsu_req_bits_ctrl_mem_unsigned,
  input  [5:0]  io_lsu_req_bits_ctrl_alu_fn,
  input         io_lsu_req_bits_ctrl_mem,
  input  [1:0]  io_lsu_req_bits_ctrl_mem_cmd,
  input  [1:0]  io_lsu_req_bits_ctrl_mop,
  input  [4:0]  io_lsu_req_bits_ctrl_reg_idxw,
  input         io_lsu_req_bits_ctrl_wfd,
  input         io_lsu_req_bits_ctrl_fence,
  input         io_lsu_req_bits_ctrl_sfu,
  input         io_lsu_req_bits_ctrl_readmask,
  input         io_lsu_req_bits_ctrl_writemask,
  input         io_lsu_req_bits_ctrl_wxd,
  input  [31:0] io_lsu_req_bits_ctrl_pc,
  output        io_dcache_rsp_ready,
  input         io_dcache_rsp_valid,
  input  [1:0]  io_dcache_rsp_bits_instrId,
  input  [31:0] io_dcache_rsp_bits_data_0,
  input  [31:0] io_dcache_rsp_bits_data_1,
  input  [31:0] io_dcache_rsp_bits_data_2,
  input  [31:0] io_dcache_rsp_bits_data_3,
  input  [31:0] io_dcache_rsp_bits_data_4,
  input  [31:0] io_dcache_rsp_bits_data_5,
  input  [31:0] io_dcache_rsp_bits_data_6,
  input  [31:0] io_dcache_rsp_bits_data_7,
  input         io_dcache_rsp_bits_activeMask_0,
  input         io_dcache_rsp_bits_activeMask_1,
  input         io_dcache_rsp_bits_activeMask_2,
  input         io_dcache_rsp_bits_activeMask_3,
  input         io_dcache_rsp_bits_activeMask_4,
  input         io_dcache_rsp_bits_activeMask_5,
  input         io_dcache_rsp_bits_activeMask_6,
  input         io_dcache_rsp_bits_activeMask_7,
  input         io_lsu_rsp_ready,
  output        io_lsu_rsp_valid,
  output [1:0]  io_lsu_rsp_bits_tag_warp_id,
  output        io_lsu_rsp_bits_tag_wfd,
  output        io_lsu_rsp_bits_tag_wxd,
  output [4:0]  io_lsu_rsp_bits_tag_reg_idxw,
  output        io_lsu_rsp_bits_tag_mask_0,
  output        io_lsu_rsp_bits_tag_mask_1,
  output        io_lsu_rsp_bits_tag_mask_2,
  output        io_lsu_rsp_bits_tag_mask_3,
  output        io_lsu_rsp_bits_tag_mask_4,
  output        io_lsu_rsp_bits_tag_mask_5,
  output        io_lsu_rsp_bits_tag_mask_6,
  output        io_lsu_rsp_bits_tag_mask_7,
  output        io_lsu_rsp_bits_tag_isWrite,
  output [31:0] io_lsu_rsp_bits_data_0,
  output [31:0] io_lsu_rsp_bits_data_1,
  output [31:0] io_lsu_rsp_bits_data_2,
  output [31:0] io_lsu_rsp_bits_data_3,
  output [31:0] io_lsu_rsp_bits_data_4,
  output [31:0] io_lsu_rsp_bits_data_5,
  output [31:0] io_lsu_rsp_bits_data_6,
  output [31:0] io_lsu_rsp_bits_data_7,
  input         io_dcache_req_ready,
  output        io_dcache_req_valid,
  output [1:0]  io_dcache_req_bits_instrId,
  output        io_dcache_req_bits_isWrite,
  output [21:0] io_dcache_req_bits_tag,
  output [4:0]  io_dcache_req_bits_setIdx,
  output        io_dcache_req_bits_perLaneAddr_0_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_0_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_1_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_1_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_2_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_2_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_3_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_3_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_4_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_4_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_5_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_5_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_6_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_6_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_7_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_7_blockOffset,
  output [31:0] io_dcache_req_bits_data_0,
  output [31:0] io_dcache_req_bits_data_1,
  output [31:0] io_dcache_req_bits_data_2,
  output [31:0] io_dcache_req_bits_data_3,
  output [31:0] io_dcache_req_bits_data_4,
  output [31:0] io_dcache_req_bits_data_5,
  output [31:0] io_dcache_req_bits_data_6,
  output [31:0] io_dcache_req_bits_data_7,
  input         io_shared_req_ready,
  output        io_shared_req_valid,
  output [1:0]  io_shared_req_bits_instrId,
  output        io_shared_req_bits_isWrite,
  output [4:0]  io_shared_req_bits_setIdx,
  output        io_shared_req_bits_perLaneAddr_0_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_0_blockOffset,
  output        io_shared_req_bits_perLaneAddr_1_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_1_blockOffset,
  output        io_shared_req_bits_perLaneAddr_2_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_2_blockOffset,
  output        io_shared_req_bits_perLaneAddr_3_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_3_blockOffset,
  output        io_shared_req_bits_perLaneAddr_4_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_4_blockOffset,
  output        io_shared_req_bits_perLaneAddr_5_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_5_blockOffset,
  output        io_shared_req_bits_perLaneAddr_6_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_6_blockOffset,
  output        io_shared_req_bits_perLaneAddr_7_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_7_blockOffset,
  output [31:0] io_shared_req_bits_data_0,
  output [31:0] io_shared_req_bits_data_1,
  output [31:0] io_shared_req_bits_data_2,
  output [31:0] io_shared_req_bits_data_3,
  output [31:0] io_shared_req_bits_data_4,
  output [31:0] io_shared_req_bits_data_5,
  output [31:0] io_shared_req_bits_data_6,
  output [31:0] io_shared_req_bits_data_7,
  output        io_shared_rsp_ready,
  input         io_shared_rsp_valid,
  input  [1:0]  io_shared_rsp_bits_instrId,
  input  [31:0] io_shared_rsp_bits_data_0,
  input  [31:0] io_shared_rsp_bits_data_1,
  input  [31:0] io_shared_rsp_bits_data_2,
  input  [31:0] io_shared_rsp_bits_data_3,
  input  [31:0] io_shared_rsp_bits_data_4,
  input  [31:0] io_shared_rsp_bits_data_5,
  input  [31:0] io_shared_rsp_bits_data_6,
  input  [31:0] io_shared_rsp_bits_data_7,
  input         io_shared_rsp_bits_activeMask_0,
  input         io_shared_rsp_bits_activeMask_1,
  input         io_shared_rsp_bits_activeMask_2,
  input         io_shared_rsp_bits_activeMask_3,
  input         io_shared_rsp_bits_activeMask_4,
  input         io_shared_rsp_bits_activeMask_5,
  input         io_shared_rsp_bits_activeMask_6,
  input         io_shared_rsp_bits_activeMask_7,
  output [3:0]  io_fence_end
);
  wire  InputFIFO_clock; // @[LSU.scala 336:25]
  wire  InputFIFO_reset; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_ready; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_valid; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_0; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_1; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_2; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_3; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_4; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_5; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_6; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in1_7; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_0; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_1; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_2; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_3; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_4; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_5; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_6; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in2_7; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_0; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_1; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_2; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_3; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_4; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_5; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_6; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_in3_7; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_0; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_1; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_2; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_3; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_4; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_5; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_6; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_mask_7; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_ctrl_inst; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_enq_bits_ctrl_wid; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_fp; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_enq_bits_ctrl_branch; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_simt_stack; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_simt_stack_op; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_barrier; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_enq_bits_ctrl_csr; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_reverse; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_isvec; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_mem_unsigned; // @[LSU.scala 336:25]
  wire [5:0] InputFIFO_io_enq_bits_ctrl_alu_fn; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_mem; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_enq_bits_ctrl_mem_cmd; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_enq_bits_ctrl_mop; // @[LSU.scala 336:25]
  wire [4:0] InputFIFO_io_enq_bits_ctrl_reg_idxw; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_wfd; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_fence; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_sfu; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_readmask; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_writemask; // @[LSU.scala 336:25]
  wire  InputFIFO_io_enq_bits_ctrl_wxd; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_enq_bits_ctrl_pc; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_ready; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_valid; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_0; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_1; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_2; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_3; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_4; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_5; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_6; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in1_7; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_0; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_1; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_2; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_3; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_4; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_5; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_6; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in2_7; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_0; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_1; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_2; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_3; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_4; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_5; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_6; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_in3_7; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_0; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_1; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_2; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_3; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_4; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_5; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_6; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_mask_7; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_ctrl_inst; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_deq_bits_ctrl_wid; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_fp; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_deq_bits_ctrl_branch; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_simt_stack; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_simt_stack_op; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_barrier; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_deq_bits_ctrl_csr; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_reverse; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_isvec; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_mem_unsigned; // @[LSU.scala 336:25]
  wire [5:0] InputFIFO_io_deq_bits_ctrl_alu_fn; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_mem; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_deq_bits_ctrl_mem_cmd; // @[LSU.scala 336:25]
  wire [1:0] InputFIFO_io_deq_bits_ctrl_mop; // @[LSU.scala 336:25]
  wire [4:0] InputFIFO_io_deq_bits_ctrl_reg_idxw; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_wfd; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_fence; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_sfu; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_readmask; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_writemask; // @[LSU.scala 336:25]
  wire  InputFIFO_io_deq_bits_ctrl_wxd; // @[LSU.scala 336:25]
  wire [31:0] InputFIFO_io_deq_bits_ctrl_pc; // @[LSU.scala 336:25]
  wire  AddrCalc_clock; // @[LSU.scala 339:24]
  wire  AddrCalc_reset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_ready; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_valid; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_0; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_1; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_2; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_3; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_4; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_5; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_6; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in1_7; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_0; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_1; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_2; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_3; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_4; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_5; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_6; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in2_7; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_0; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_1; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_2; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_3; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_4; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_5; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_6; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_from_fifo_bits_in3_7; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_0; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_1; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_2; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_3; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_4; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_5; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_6; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_mask_7; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_from_fifo_bits_ctrl_wid; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_ctrl_isvec; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_ctrl_mem_unsigned; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_from_fifo_bits_ctrl_mem_cmd; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_from_fifo_bits_ctrl_mop; // @[LSU.scala 339:24]
  wire [4:0] AddrCalc_io_from_fifo_bits_ctrl_reg_idxw; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_ctrl_wfd; // @[LSU.scala 339:24]
  wire  AddrCalc_io_from_fifo_bits_ctrl_wxd; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_ready; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_valid; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_to_mshr_bits_tag_warp_id; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_wfd; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_wxd; // @[LSU.scala 339:24]
  wire [4:0] AddrCalc_io_to_mshr_bits_tag_reg_idxw; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_0; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_1; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_2; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_3; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_4; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_5; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_6; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_mask_7; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_unsigned; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_isvec; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_mshr_bits_tag_isWrite; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_idx_entry; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_ready; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_valid; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_to_dcache_bits_instrId; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_isWrite; // @[LSU.scala 339:24]
  wire [21:0] AddrCalc_io_to_dcache_bits_tag; // @[LSU.scala 339:24]
  wire [4:0] AddrCalc_io_to_dcache_bits_setIdx; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_0_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_0_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_1_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_1_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_2_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_2_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_3_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_3_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_4_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_4_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_5_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_5_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_6_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_6_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_dcache_bits_perLaneAddr_7_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_dcache_bits_perLaneAddr_7_blockOffset; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_0; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_1; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_2; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_3; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_4; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_5; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_6; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_dcache_bits_data_7; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_ready; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_valid; // @[LSU.scala 339:24]
  wire [1:0] AddrCalc_io_to_shared_bits_instrId; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_isWrite; // @[LSU.scala 339:24]
  wire [4:0] AddrCalc_io_to_shared_bits_setIdx; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_0_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_0_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_1_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_1_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_2_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_2_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_3_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_3_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_4_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_4_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_5_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_5_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_6_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_6_blockOffset; // @[LSU.scala 339:24]
  wire  AddrCalc_io_to_shared_bits_perLaneAddr_7_activeMask; // @[LSU.scala 339:24]
  wire [2:0] AddrCalc_io_to_shared_bits_perLaneAddr_7_blockOffset; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_0; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_1; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_2; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_3; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_4; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_5; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_6; // @[LSU.scala 339:24]
  wire [31:0] AddrCalc_io_to_shared_bits_data_7; // @[LSU.scala 339:24]
  wire  rspArbiter_io_in_0_ready; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_valid; // @[LSU.scala 344:26]
  wire [1:0] rspArbiter_io_in_0_bits_instrId; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_0; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_1; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_2; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_3; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_4; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_5; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_6; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_0_bits_data_7; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_0; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_1; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_2; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_3; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_4; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_5; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_6; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_0_bits_activeMask_7; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_ready; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_valid; // @[LSU.scala 344:26]
  wire [1:0] rspArbiter_io_in_1_bits_instrId; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_0; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_1; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_2; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_3; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_4; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_5; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_6; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_in_1_bits_data_7; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_0; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_1; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_2; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_3; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_4; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_5; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_6; // @[LSU.scala 344:26]
  wire  rspArbiter_io_in_1_bits_activeMask_7; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_ready; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_valid; // @[LSU.scala 344:26]
  wire [1:0] rspArbiter_io_out_bits_instrId; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_0; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_1; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_2; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_3; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_4; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_5; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_6; // @[LSU.scala 344:26]
  wire [31:0] rspArbiter_io_out_bits_data_7; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_0; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_1; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_2; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_3; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_4; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_5; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_6; // @[LSU.scala 344:26]
  wire  rspArbiter_io_out_bits_activeMask_7; // @[LSU.scala 344:26]
  wire  Coalscer_clock; // @[LSU.scala 349:24]
  wire  Coalscer_reset; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_ready; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_valid; // @[LSU.scala 349:24]
  wire [1:0] Coalscer_io_from_addr_bits_tag_warp_id; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_wfd; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_wxd; // @[LSU.scala 349:24]
  wire [4:0] Coalscer_io_from_addr_bits_tag_reg_idxw; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_0; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_1; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_2; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_3; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_4; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_5; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_6; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_mask_7; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_unsigned; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_isvec; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_addr_bits_tag_isWrite; // @[LSU.scala 349:24]
  wire [1:0] Coalscer_io_idx_entry; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_ready; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_valid; // @[LSU.scala 349:24]
  wire [1:0] Coalscer_io_from_dcache_bits_instrId; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_0; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_1; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_2; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_3; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_4; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_5; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_6; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_from_dcache_bits_data_7; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_0; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_1; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_2; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_3; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_4; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_5; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_6; // @[LSU.scala 349:24]
  wire  Coalscer_io_from_dcache_bits_activeMask_7; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_ready; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_valid; // @[LSU.scala 349:24]
  wire [1:0] Coalscer_io_to_pipe_bits_tag_warp_id; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_wfd; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_wxd; // @[LSU.scala 349:24]
  wire [4:0] Coalscer_io_to_pipe_bits_tag_reg_idxw; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_0; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_1; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_2; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_3; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_4; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_5; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_6; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_mask_7; // @[LSU.scala 349:24]
  wire  Coalscer_io_to_pipe_bits_tag_isWrite; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_0; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_1; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_2; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_3; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_4; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_5; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_6; // @[LSU.scala 349:24]
  wire [31:0] Coalscer_io_to_pipe_bits_data_7; // @[LSU.scala 349:24]
  wire  ShiftBoard_clock; // @[LSU.scala 356:51]
  wire  ShiftBoard_reset; // @[LSU.scala 356:51]
  wire  ShiftBoard_io_left; // @[LSU.scala 356:51]
  wire  ShiftBoard_io_right; // @[LSU.scala 356:51]
  wire  ShiftBoard_io_full; // @[LSU.scala 356:51]
  wire  ShiftBoard_io_empty; // @[LSU.scala 356:51]
  wire  ShiftBoard_1_clock; // @[LSU.scala 356:51]
  wire  ShiftBoard_1_reset; // @[LSU.scala 356:51]
  wire  ShiftBoard_1_io_left; // @[LSU.scala 356:51]
  wire  ShiftBoard_1_io_right; // @[LSU.scala 356:51]
  wire  ShiftBoard_1_io_full; // @[LSU.scala 356:51]
  wire  ShiftBoard_1_io_empty; // @[LSU.scala 356:51]
  wire  ShiftBoard_2_clock; // @[LSU.scala 356:51]
  wire  ShiftBoard_2_reset; // @[LSU.scala 356:51]
  wire  ShiftBoard_2_io_left; // @[LSU.scala 356:51]
  wire  ShiftBoard_2_io_right; // @[LSU.scala 356:51]
  wire  ShiftBoard_2_io_full; // @[LSU.scala 356:51]
  wire  ShiftBoard_2_io_empty; // @[LSU.scala 356:51]
  wire  ShiftBoard_3_clock; // @[LSU.scala 356:51]
  wire  ShiftBoard_3_reset; // @[LSU.scala 356:51]
  wire  ShiftBoard_3_io_left; // @[LSU.scala 356:51]
  wire  ShiftBoard_3_io_right; // @[LSU.scala 356:51]
  wire  ShiftBoard_3_io_full; // @[LSU.scala 356:51]
  wire  ShiftBoard_3_io_empty; // @[LSU.scala 356:51]
  wire  _shiftBoard_0_left_T = io_lsu_req_ready & io_lsu_req_valid; // @[Decoupled.scala 50:35]
  wire  _shiftBoard_0_right_T = io_lsu_rsp_ready & io_lsu_rsp_valid; // @[Decoupled.scala 50:35]
  wire  shiftBoard_1_empty = ShiftBoard_1_io_empty; // @[LSU.scala 356:{25,25}]
  wire  shiftBoard_0_empty = ShiftBoard_io_empty; // @[LSU.scala 356:{25,25}]
  wire [1:0] io_fence_end_lo = {shiftBoard_1_empty,shiftBoard_0_empty}; // @[LSU.scala 361:59]
  wire  shiftBoard_3_empty = ShiftBoard_3_io_empty; // @[LSU.scala 356:{25,25}]
  wire  shiftBoard_2_empty = ShiftBoard_2_io_empty; // @[LSU.scala 356:{25,25}]
  wire [1:0] io_fence_end_hi = {shiftBoard_3_empty,shiftBoard_2_empty}; // @[LSU.scala 361:59]
  wire  shiftBoard_0_full = ShiftBoard_io_full; // @[LSU.scala 356:{25,25}]
  wire  shiftBoard_1_full = ShiftBoard_1_io_full; // @[LSU.scala 356:{25,25}]
  wire  _GEN_1 = 2'h1 == io_lsu_req_bits_ctrl_wid ? shiftBoard_1_full : shiftBoard_0_full; // @[LSU.scala 362:{24,24}]
  wire  shiftBoard_2_full = ShiftBoard_2_io_full; // @[LSU.scala 356:{25,25}]
  wire  _GEN_2 = 2'h2 == io_lsu_req_bits_ctrl_wid ? shiftBoard_2_full : _GEN_1; // @[LSU.scala 362:{24,24}]
  wire  shiftBoard_3_full = ShiftBoard_3_io_full; // @[LSU.scala 356:{25,25}]
  wire  _GEN_3 = 2'h3 == io_lsu_req_bits_ctrl_wid ? shiftBoard_3_full : _GEN_2; // @[LSU.scala 362:{24,24}]
  Queue_41 InputFIFO ( // @[LSU.scala 336:25]
    .clock(InputFIFO_clock),
    .reset(InputFIFO_reset),
    .io_enq_ready(InputFIFO_io_enq_ready),
    .io_enq_valid(InputFIFO_io_enq_valid),
    .io_enq_bits_in1_0(InputFIFO_io_enq_bits_in1_0),
    .io_enq_bits_in1_1(InputFIFO_io_enq_bits_in1_1),
    .io_enq_bits_in1_2(InputFIFO_io_enq_bits_in1_2),
    .io_enq_bits_in1_3(InputFIFO_io_enq_bits_in1_3),
    .io_enq_bits_in1_4(InputFIFO_io_enq_bits_in1_4),
    .io_enq_bits_in1_5(InputFIFO_io_enq_bits_in1_5),
    .io_enq_bits_in1_6(InputFIFO_io_enq_bits_in1_6),
    .io_enq_bits_in1_7(InputFIFO_io_enq_bits_in1_7),
    .io_enq_bits_in2_0(InputFIFO_io_enq_bits_in2_0),
    .io_enq_bits_in2_1(InputFIFO_io_enq_bits_in2_1),
    .io_enq_bits_in2_2(InputFIFO_io_enq_bits_in2_2),
    .io_enq_bits_in2_3(InputFIFO_io_enq_bits_in2_3),
    .io_enq_bits_in2_4(InputFIFO_io_enq_bits_in2_4),
    .io_enq_bits_in2_5(InputFIFO_io_enq_bits_in2_5),
    .io_enq_bits_in2_6(InputFIFO_io_enq_bits_in2_6),
    .io_enq_bits_in2_7(InputFIFO_io_enq_bits_in2_7),
    .io_enq_bits_in3_0(InputFIFO_io_enq_bits_in3_0),
    .io_enq_bits_in3_1(InputFIFO_io_enq_bits_in3_1),
    .io_enq_bits_in3_2(InputFIFO_io_enq_bits_in3_2),
    .io_enq_bits_in3_3(InputFIFO_io_enq_bits_in3_3),
    .io_enq_bits_in3_4(InputFIFO_io_enq_bits_in3_4),
    .io_enq_bits_in3_5(InputFIFO_io_enq_bits_in3_5),
    .io_enq_bits_in3_6(InputFIFO_io_enq_bits_in3_6),
    .io_enq_bits_in3_7(InputFIFO_io_enq_bits_in3_7),
    .io_enq_bits_mask_0(InputFIFO_io_enq_bits_mask_0),
    .io_enq_bits_mask_1(InputFIFO_io_enq_bits_mask_1),
    .io_enq_bits_mask_2(InputFIFO_io_enq_bits_mask_2),
    .io_enq_bits_mask_3(InputFIFO_io_enq_bits_mask_3),
    .io_enq_bits_mask_4(InputFIFO_io_enq_bits_mask_4),
    .io_enq_bits_mask_5(InputFIFO_io_enq_bits_mask_5),
    .io_enq_bits_mask_6(InputFIFO_io_enq_bits_mask_6),
    .io_enq_bits_mask_7(InputFIFO_io_enq_bits_mask_7),
    .io_enq_bits_ctrl_inst(InputFIFO_io_enq_bits_ctrl_inst),
    .io_enq_bits_ctrl_wid(InputFIFO_io_enq_bits_ctrl_wid),
    .io_enq_bits_ctrl_fp(InputFIFO_io_enq_bits_ctrl_fp),
    .io_enq_bits_ctrl_branch(InputFIFO_io_enq_bits_ctrl_branch),
    .io_enq_bits_ctrl_simt_stack(InputFIFO_io_enq_bits_ctrl_simt_stack),
    .io_enq_bits_ctrl_simt_stack_op(InputFIFO_io_enq_bits_ctrl_simt_stack_op),
    .io_enq_bits_ctrl_barrier(InputFIFO_io_enq_bits_ctrl_barrier),
    .io_enq_bits_ctrl_csr(InputFIFO_io_enq_bits_ctrl_csr),
    .io_enq_bits_ctrl_reverse(InputFIFO_io_enq_bits_ctrl_reverse),
    .io_enq_bits_ctrl_isvec(InputFIFO_io_enq_bits_ctrl_isvec),
    .io_enq_bits_ctrl_mem_unsigned(InputFIFO_io_enq_bits_ctrl_mem_unsigned),
    .io_enq_bits_ctrl_alu_fn(InputFIFO_io_enq_bits_ctrl_alu_fn),
    .io_enq_bits_ctrl_mem(InputFIFO_io_enq_bits_ctrl_mem),
    .io_enq_bits_ctrl_mem_cmd(InputFIFO_io_enq_bits_ctrl_mem_cmd),
    .io_enq_bits_ctrl_mop(InputFIFO_io_enq_bits_ctrl_mop),
    .io_enq_bits_ctrl_reg_idxw(InputFIFO_io_enq_bits_ctrl_reg_idxw),
    .io_enq_bits_ctrl_wfd(InputFIFO_io_enq_bits_ctrl_wfd),
    .io_enq_bits_ctrl_fence(InputFIFO_io_enq_bits_ctrl_fence),
    .io_enq_bits_ctrl_sfu(InputFIFO_io_enq_bits_ctrl_sfu),
    .io_enq_bits_ctrl_readmask(InputFIFO_io_enq_bits_ctrl_readmask),
    .io_enq_bits_ctrl_writemask(InputFIFO_io_enq_bits_ctrl_writemask),
    .io_enq_bits_ctrl_wxd(InputFIFO_io_enq_bits_ctrl_wxd),
    .io_enq_bits_ctrl_pc(InputFIFO_io_enq_bits_ctrl_pc),
    .io_deq_ready(InputFIFO_io_deq_ready),
    .io_deq_valid(InputFIFO_io_deq_valid),
    .io_deq_bits_in1_0(InputFIFO_io_deq_bits_in1_0),
    .io_deq_bits_in1_1(InputFIFO_io_deq_bits_in1_1),
    .io_deq_bits_in1_2(InputFIFO_io_deq_bits_in1_2),
    .io_deq_bits_in1_3(InputFIFO_io_deq_bits_in1_3),
    .io_deq_bits_in1_4(InputFIFO_io_deq_bits_in1_4),
    .io_deq_bits_in1_5(InputFIFO_io_deq_bits_in1_5),
    .io_deq_bits_in1_6(InputFIFO_io_deq_bits_in1_6),
    .io_deq_bits_in1_7(InputFIFO_io_deq_bits_in1_7),
    .io_deq_bits_in2_0(InputFIFO_io_deq_bits_in2_0),
    .io_deq_bits_in2_1(InputFIFO_io_deq_bits_in2_1),
    .io_deq_bits_in2_2(InputFIFO_io_deq_bits_in2_2),
    .io_deq_bits_in2_3(InputFIFO_io_deq_bits_in2_3),
    .io_deq_bits_in2_4(InputFIFO_io_deq_bits_in2_4),
    .io_deq_bits_in2_5(InputFIFO_io_deq_bits_in2_5),
    .io_deq_bits_in2_6(InputFIFO_io_deq_bits_in2_6),
    .io_deq_bits_in2_7(InputFIFO_io_deq_bits_in2_7),
    .io_deq_bits_in3_0(InputFIFO_io_deq_bits_in3_0),
    .io_deq_bits_in3_1(InputFIFO_io_deq_bits_in3_1),
    .io_deq_bits_in3_2(InputFIFO_io_deq_bits_in3_2),
    .io_deq_bits_in3_3(InputFIFO_io_deq_bits_in3_3),
    .io_deq_bits_in3_4(InputFIFO_io_deq_bits_in3_4),
    .io_deq_bits_in3_5(InputFIFO_io_deq_bits_in3_5),
    .io_deq_bits_in3_6(InputFIFO_io_deq_bits_in3_6),
    .io_deq_bits_in3_7(InputFIFO_io_deq_bits_in3_7),
    .io_deq_bits_mask_0(InputFIFO_io_deq_bits_mask_0),
    .io_deq_bits_mask_1(InputFIFO_io_deq_bits_mask_1),
    .io_deq_bits_mask_2(InputFIFO_io_deq_bits_mask_2),
    .io_deq_bits_mask_3(InputFIFO_io_deq_bits_mask_3),
    .io_deq_bits_mask_4(InputFIFO_io_deq_bits_mask_4),
    .io_deq_bits_mask_5(InputFIFO_io_deq_bits_mask_5),
    .io_deq_bits_mask_6(InputFIFO_io_deq_bits_mask_6),
    .io_deq_bits_mask_7(InputFIFO_io_deq_bits_mask_7),
    .io_deq_bits_ctrl_inst(InputFIFO_io_deq_bits_ctrl_inst),
    .io_deq_bits_ctrl_wid(InputFIFO_io_deq_bits_ctrl_wid),
    .io_deq_bits_ctrl_fp(InputFIFO_io_deq_bits_ctrl_fp),
    .io_deq_bits_ctrl_branch(InputFIFO_io_deq_bits_ctrl_branch),
    .io_deq_bits_ctrl_simt_stack(InputFIFO_io_deq_bits_ctrl_simt_stack),
    .io_deq_bits_ctrl_simt_stack_op(InputFIFO_io_deq_bits_ctrl_simt_stack_op),
    .io_deq_bits_ctrl_barrier(InputFIFO_io_deq_bits_ctrl_barrier),
    .io_deq_bits_ctrl_csr(InputFIFO_io_deq_bits_ctrl_csr),
    .io_deq_bits_ctrl_reverse(InputFIFO_io_deq_bits_ctrl_reverse),
    .io_deq_bits_ctrl_isvec(InputFIFO_io_deq_bits_ctrl_isvec),
    .io_deq_bits_ctrl_mem_unsigned(InputFIFO_io_deq_bits_ctrl_mem_unsigned),
    .io_deq_bits_ctrl_alu_fn(InputFIFO_io_deq_bits_ctrl_alu_fn),
    .io_deq_bits_ctrl_mem(InputFIFO_io_deq_bits_ctrl_mem),
    .io_deq_bits_ctrl_mem_cmd(InputFIFO_io_deq_bits_ctrl_mem_cmd),
    .io_deq_bits_ctrl_mop(InputFIFO_io_deq_bits_ctrl_mop),
    .io_deq_bits_ctrl_reg_idxw(InputFIFO_io_deq_bits_ctrl_reg_idxw),
    .io_deq_bits_ctrl_wfd(InputFIFO_io_deq_bits_ctrl_wfd),
    .io_deq_bits_ctrl_fence(InputFIFO_io_deq_bits_ctrl_fence),
    .io_deq_bits_ctrl_sfu(InputFIFO_io_deq_bits_ctrl_sfu),
    .io_deq_bits_ctrl_readmask(InputFIFO_io_deq_bits_ctrl_readmask),
    .io_deq_bits_ctrl_writemask(InputFIFO_io_deq_bits_ctrl_writemask),
    .io_deq_bits_ctrl_wxd(InputFIFO_io_deq_bits_ctrl_wxd),
    .io_deq_bits_ctrl_pc(InputFIFO_io_deq_bits_ctrl_pc)
  );
  AddrCalculate AddrCalc ( // @[LSU.scala 339:24]
    .clock(AddrCalc_clock),
    .reset(AddrCalc_reset),
    .io_from_fifo_ready(AddrCalc_io_from_fifo_ready),
    .io_from_fifo_valid(AddrCalc_io_from_fifo_valid),
    .io_from_fifo_bits_in1_0(AddrCalc_io_from_fifo_bits_in1_0),
    .io_from_fifo_bits_in1_1(AddrCalc_io_from_fifo_bits_in1_1),
    .io_from_fifo_bits_in1_2(AddrCalc_io_from_fifo_bits_in1_2),
    .io_from_fifo_bits_in1_3(AddrCalc_io_from_fifo_bits_in1_3),
    .io_from_fifo_bits_in1_4(AddrCalc_io_from_fifo_bits_in1_4),
    .io_from_fifo_bits_in1_5(AddrCalc_io_from_fifo_bits_in1_5),
    .io_from_fifo_bits_in1_6(AddrCalc_io_from_fifo_bits_in1_6),
    .io_from_fifo_bits_in1_7(AddrCalc_io_from_fifo_bits_in1_7),
    .io_from_fifo_bits_in2_0(AddrCalc_io_from_fifo_bits_in2_0),
    .io_from_fifo_bits_in2_1(AddrCalc_io_from_fifo_bits_in2_1),
    .io_from_fifo_bits_in2_2(AddrCalc_io_from_fifo_bits_in2_2),
    .io_from_fifo_bits_in2_3(AddrCalc_io_from_fifo_bits_in2_3),
    .io_from_fifo_bits_in2_4(AddrCalc_io_from_fifo_bits_in2_4),
    .io_from_fifo_bits_in2_5(AddrCalc_io_from_fifo_bits_in2_5),
    .io_from_fifo_bits_in2_6(AddrCalc_io_from_fifo_bits_in2_6),
    .io_from_fifo_bits_in2_7(AddrCalc_io_from_fifo_bits_in2_7),
    .io_from_fifo_bits_in3_0(AddrCalc_io_from_fifo_bits_in3_0),
    .io_from_fifo_bits_in3_1(AddrCalc_io_from_fifo_bits_in3_1),
    .io_from_fifo_bits_in3_2(AddrCalc_io_from_fifo_bits_in3_2),
    .io_from_fifo_bits_in3_3(AddrCalc_io_from_fifo_bits_in3_3),
    .io_from_fifo_bits_in3_4(AddrCalc_io_from_fifo_bits_in3_4),
    .io_from_fifo_bits_in3_5(AddrCalc_io_from_fifo_bits_in3_5),
    .io_from_fifo_bits_in3_6(AddrCalc_io_from_fifo_bits_in3_6),
    .io_from_fifo_bits_in3_7(AddrCalc_io_from_fifo_bits_in3_7),
    .io_from_fifo_bits_mask_0(AddrCalc_io_from_fifo_bits_mask_0),
    .io_from_fifo_bits_mask_1(AddrCalc_io_from_fifo_bits_mask_1),
    .io_from_fifo_bits_mask_2(AddrCalc_io_from_fifo_bits_mask_2),
    .io_from_fifo_bits_mask_3(AddrCalc_io_from_fifo_bits_mask_3),
    .io_from_fifo_bits_mask_4(AddrCalc_io_from_fifo_bits_mask_4),
    .io_from_fifo_bits_mask_5(AddrCalc_io_from_fifo_bits_mask_5),
    .io_from_fifo_bits_mask_6(AddrCalc_io_from_fifo_bits_mask_6),
    .io_from_fifo_bits_mask_7(AddrCalc_io_from_fifo_bits_mask_7),
    .io_from_fifo_bits_ctrl_wid(AddrCalc_io_from_fifo_bits_ctrl_wid),
    .io_from_fifo_bits_ctrl_isvec(AddrCalc_io_from_fifo_bits_ctrl_isvec),
    .io_from_fifo_bits_ctrl_mem_unsigned(AddrCalc_io_from_fifo_bits_ctrl_mem_unsigned),
    .io_from_fifo_bits_ctrl_mem_cmd(AddrCalc_io_from_fifo_bits_ctrl_mem_cmd),
    .io_from_fifo_bits_ctrl_mop(AddrCalc_io_from_fifo_bits_ctrl_mop),
    .io_from_fifo_bits_ctrl_reg_idxw(AddrCalc_io_from_fifo_bits_ctrl_reg_idxw),
    .io_from_fifo_bits_ctrl_wfd(AddrCalc_io_from_fifo_bits_ctrl_wfd),
    .io_from_fifo_bits_ctrl_wxd(AddrCalc_io_from_fifo_bits_ctrl_wxd),
    .io_to_mshr_ready(AddrCalc_io_to_mshr_ready),
    .io_to_mshr_valid(AddrCalc_io_to_mshr_valid),
    .io_to_mshr_bits_tag_warp_id(AddrCalc_io_to_mshr_bits_tag_warp_id),
    .io_to_mshr_bits_tag_wfd(AddrCalc_io_to_mshr_bits_tag_wfd),
    .io_to_mshr_bits_tag_wxd(AddrCalc_io_to_mshr_bits_tag_wxd),
    .io_to_mshr_bits_tag_reg_idxw(AddrCalc_io_to_mshr_bits_tag_reg_idxw),
    .io_to_mshr_bits_tag_mask_0(AddrCalc_io_to_mshr_bits_tag_mask_0),
    .io_to_mshr_bits_tag_mask_1(AddrCalc_io_to_mshr_bits_tag_mask_1),
    .io_to_mshr_bits_tag_mask_2(AddrCalc_io_to_mshr_bits_tag_mask_2),
    .io_to_mshr_bits_tag_mask_3(AddrCalc_io_to_mshr_bits_tag_mask_3),
    .io_to_mshr_bits_tag_mask_4(AddrCalc_io_to_mshr_bits_tag_mask_4),
    .io_to_mshr_bits_tag_mask_5(AddrCalc_io_to_mshr_bits_tag_mask_5),
    .io_to_mshr_bits_tag_mask_6(AddrCalc_io_to_mshr_bits_tag_mask_6),
    .io_to_mshr_bits_tag_mask_7(AddrCalc_io_to_mshr_bits_tag_mask_7),
    .io_to_mshr_bits_tag_unsigned(AddrCalc_io_to_mshr_bits_tag_unsigned),
    .io_to_mshr_bits_tag_isvec(AddrCalc_io_to_mshr_bits_tag_isvec),
    .io_to_mshr_bits_tag_isWrite(AddrCalc_io_to_mshr_bits_tag_isWrite),
    .io_idx_entry(AddrCalc_io_idx_entry),
    .io_to_dcache_ready(AddrCalc_io_to_dcache_ready),
    .io_to_dcache_valid(AddrCalc_io_to_dcache_valid),
    .io_to_dcache_bits_instrId(AddrCalc_io_to_dcache_bits_instrId),
    .io_to_dcache_bits_isWrite(AddrCalc_io_to_dcache_bits_isWrite),
    .io_to_dcache_bits_tag(AddrCalc_io_to_dcache_bits_tag),
    .io_to_dcache_bits_setIdx(AddrCalc_io_to_dcache_bits_setIdx),
    .io_to_dcache_bits_perLaneAddr_0_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_0_activeMask),
    .io_to_dcache_bits_perLaneAddr_0_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_0_blockOffset),
    .io_to_dcache_bits_perLaneAddr_1_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_1_activeMask),
    .io_to_dcache_bits_perLaneAddr_1_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_1_blockOffset),
    .io_to_dcache_bits_perLaneAddr_2_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_2_activeMask),
    .io_to_dcache_bits_perLaneAddr_2_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_2_blockOffset),
    .io_to_dcache_bits_perLaneAddr_3_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_3_activeMask),
    .io_to_dcache_bits_perLaneAddr_3_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_3_blockOffset),
    .io_to_dcache_bits_perLaneAddr_4_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_4_activeMask),
    .io_to_dcache_bits_perLaneAddr_4_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_4_blockOffset),
    .io_to_dcache_bits_perLaneAddr_5_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_5_activeMask),
    .io_to_dcache_bits_perLaneAddr_5_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_5_blockOffset),
    .io_to_dcache_bits_perLaneAddr_6_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_6_activeMask),
    .io_to_dcache_bits_perLaneAddr_6_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_6_blockOffset),
    .io_to_dcache_bits_perLaneAddr_7_activeMask(AddrCalc_io_to_dcache_bits_perLaneAddr_7_activeMask),
    .io_to_dcache_bits_perLaneAddr_7_blockOffset(AddrCalc_io_to_dcache_bits_perLaneAddr_7_blockOffset),
    .io_to_dcache_bits_data_0(AddrCalc_io_to_dcache_bits_data_0),
    .io_to_dcache_bits_data_1(AddrCalc_io_to_dcache_bits_data_1),
    .io_to_dcache_bits_data_2(AddrCalc_io_to_dcache_bits_data_2),
    .io_to_dcache_bits_data_3(AddrCalc_io_to_dcache_bits_data_3),
    .io_to_dcache_bits_data_4(AddrCalc_io_to_dcache_bits_data_4),
    .io_to_dcache_bits_data_5(AddrCalc_io_to_dcache_bits_data_5),
    .io_to_dcache_bits_data_6(AddrCalc_io_to_dcache_bits_data_6),
    .io_to_dcache_bits_data_7(AddrCalc_io_to_dcache_bits_data_7),
    .io_to_shared_ready(AddrCalc_io_to_shared_ready),
    .io_to_shared_valid(AddrCalc_io_to_shared_valid),
    .io_to_shared_bits_instrId(AddrCalc_io_to_shared_bits_instrId),
    .io_to_shared_bits_isWrite(AddrCalc_io_to_shared_bits_isWrite),
    .io_to_shared_bits_setIdx(AddrCalc_io_to_shared_bits_setIdx),
    .io_to_shared_bits_perLaneAddr_0_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_0_activeMask),
    .io_to_shared_bits_perLaneAddr_0_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_0_blockOffset),
    .io_to_shared_bits_perLaneAddr_1_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_1_activeMask),
    .io_to_shared_bits_perLaneAddr_1_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_1_blockOffset),
    .io_to_shared_bits_perLaneAddr_2_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_2_activeMask),
    .io_to_shared_bits_perLaneAddr_2_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_2_blockOffset),
    .io_to_shared_bits_perLaneAddr_3_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_3_activeMask),
    .io_to_shared_bits_perLaneAddr_3_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_3_blockOffset),
    .io_to_shared_bits_perLaneAddr_4_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_4_activeMask),
    .io_to_shared_bits_perLaneAddr_4_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_4_blockOffset),
    .io_to_shared_bits_perLaneAddr_5_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_5_activeMask),
    .io_to_shared_bits_perLaneAddr_5_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_5_blockOffset),
    .io_to_shared_bits_perLaneAddr_6_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_6_activeMask),
    .io_to_shared_bits_perLaneAddr_6_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_6_blockOffset),
    .io_to_shared_bits_perLaneAddr_7_activeMask(AddrCalc_io_to_shared_bits_perLaneAddr_7_activeMask),
    .io_to_shared_bits_perLaneAddr_7_blockOffset(AddrCalc_io_to_shared_bits_perLaneAddr_7_blockOffset),
    .io_to_shared_bits_data_0(AddrCalc_io_to_shared_bits_data_0),
    .io_to_shared_bits_data_1(AddrCalc_io_to_shared_bits_data_1),
    .io_to_shared_bits_data_2(AddrCalc_io_to_shared_bits_data_2),
    .io_to_shared_bits_data_3(AddrCalc_io_to_shared_bits_data_3),
    .io_to_shared_bits_data_4(AddrCalc_io_to_shared_bits_data_4),
    .io_to_shared_bits_data_5(AddrCalc_io_to_shared_bits_data_5),
    .io_to_shared_bits_data_6(AddrCalc_io_to_shared_bits_data_6),
    .io_to_shared_bits_data_7(AddrCalc_io_to_shared_bits_data_7)
  );
  Arbiter_8 rspArbiter ( // @[LSU.scala 344:26]
    .io_in_0_ready(rspArbiter_io_in_0_ready),
    .io_in_0_valid(rspArbiter_io_in_0_valid),
    .io_in_0_bits_instrId(rspArbiter_io_in_0_bits_instrId),
    .io_in_0_bits_data_0(rspArbiter_io_in_0_bits_data_0),
    .io_in_0_bits_data_1(rspArbiter_io_in_0_bits_data_1),
    .io_in_0_bits_data_2(rspArbiter_io_in_0_bits_data_2),
    .io_in_0_bits_data_3(rspArbiter_io_in_0_bits_data_3),
    .io_in_0_bits_data_4(rspArbiter_io_in_0_bits_data_4),
    .io_in_0_bits_data_5(rspArbiter_io_in_0_bits_data_5),
    .io_in_0_bits_data_6(rspArbiter_io_in_0_bits_data_6),
    .io_in_0_bits_data_7(rspArbiter_io_in_0_bits_data_7),
    .io_in_0_bits_activeMask_0(rspArbiter_io_in_0_bits_activeMask_0),
    .io_in_0_bits_activeMask_1(rspArbiter_io_in_0_bits_activeMask_1),
    .io_in_0_bits_activeMask_2(rspArbiter_io_in_0_bits_activeMask_2),
    .io_in_0_bits_activeMask_3(rspArbiter_io_in_0_bits_activeMask_3),
    .io_in_0_bits_activeMask_4(rspArbiter_io_in_0_bits_activeMask_4),
    .io_in_0_bits_activeMask_5(rspArbiter_io_in_0_bits_activeMask_5),
    .io_in_0_bits_activeMask_6(rspArbiter_io_in_0_bits_activeMask_6),
    .io_in_0_bits_activeMask_7(rspArbiter_io_in_0_bits_activeMask_7),
    .io_in_1_ready(rspArbiter_io_in_1_ready),
    .io_in_1_valid(rspArbiter_io_in_1_valid),
    .io_in_1_bits_instrId(rspArbiter_io_in_1_bits_instrId),
    .io_in_1_bits_data_0(rspArbiter_io_in_1_bits_data_0),
    .io_in_1_bits_data_1(rspArbiter_io_in_1_bits_data_1),
    .io_in_1_bits_data_2(rspArbiter_io_in_1_bits_data_2),
    .io_in_1_bits_data_3(rspArbiter_io_in_1_bits_data_3),
    .io_in_1_bits_data_4(rspArbiter_io_in_1_bits_data_4),
    .io_in_1_bits_data_5(rspArbiter_io_in_1_bits_data_5),
    .io_in_1_bits_data_6(rspArbiter_io_in_1_bits_data_6),
    .io_in_1_bits_data_7(rspArbiter_io_in_1_bits_data_7),
    .io_in_1_bits_activeMask_0(rspArbiter_io_in_1_bits_activeMask_0),
    .io_in_1_bits_activeMask_1(rspArbiter_io_in_1_bits_activeMask_1),
    .io_in_1_bits_activeMask_2(rspArbiter_io_in_1_bits_activeMask_2),
    .io_in_1_bits_activeMask_3(rspArbiter_io_in_1_bits_activeMask_3),
    .io_in_1_bits_activeMask_4(rspArbiter_io_in_1_bits_activeMask_4),
    .io_in_1_bits_activeMask_5(rspArbiter_io_in_1_bits_activeMask_5),
    .io_in_1_bits_activeMask_6(rspArbiter_io_in_1_bits_activeMask_6),
    .io_in_1_bits_activeMask_7(rspArbiter_io_in_1_bits_activeMask_7),
    .io_out_ready(rspArbiter_io_out_ready),
    .io_out_valid(rspArbiter_io_out_valid),
    .io_out_bits_instrId(rspArbiter_io_out_bits_instrId),
    .io_out_bits_data_0(rspArbiter_io_out_bits_data_0),
    .io_out_bits_data_1(rspArbiter_io_out_bits_data_1),
    .io_out_bits_data_2(rspArbiter_io_out_bits_data_2),
    .io_out_bits_data_3(rspArbiter_io_out_bits_data_3),
    .io_out_bits_data_4(rspArbiter_io_out_bits_data_4),
    .io_out_bits_data_5(rspArbiter_io_out_bits_data_5),
    .io_out_bits_data_6(rspArbiter_io_out_bits_data_6),
    .io_out_bits_data_7(rspArbiter_io_out_bits_data_7),
    .io_out_bits_activeMask_0(rspArbiter_io_out_bits_activeMask_0),
    .io_out_bits_activeMask_1(rspArbiter_io_out_bits_activeMask_1),
    .io_out_bits_activeMask_2(rspArbiter_io_out_bits_activeMask_2),
    .io_out_bits_activeMask_3(rspArbiter_io_out_bits_activeMask_3),
    .io_out_bits_activeMask_4(rspArbiter_io_out_bits_activeMask_4),
    .io_out_bits_activeMask_5(rspArbiter_io_out_bits_activeMask_5),
    .io_out_bits_activeMask_6(rspArbiter_io_out_bits_activeMask_6),
    .io_out_bits_activeMask_7(rspArbiter_io_out_bits_activeMask_7)
  );
  MSHRv2 Coalscer ( // @[LSU.scala 349:24]
    .clock(Coalscer_clock),
    .reset(Coalscer_reset),
    .io_from_addr_ready(Coalscer_io_from_addr_ready),
    .io_from_addr_valid(Coalscer_io_from_addr_valid),
    .io_from_addr_bits_tag_warp_id(Coalscer_io_from_addr_bits_tag_warp_id),
    .io_from_addr_bits_tag_wfd(Coalscer_io_from_addr_bits_tag_wfd),
    .io_from_addr_bits_tag_wxd(Coalscer_io_from_addr_bits_tag_wxd),
    .io_from_addr_bits_tag_reg_idxw(Coalscer_io_from_addr_bits_tag_reg_idxw),
    .io_from_addr_bits_tag_mask_0(Coalscer_io_from_addr_bits_tag_mask_0),
    .io_from_addr_bits_tag_mask_1(Coalscer_io_from_addr_bits_tag_mask_1),
    .io_from_addr_bits_tag_mask_2(Coalscer_io_from_addr_bits_tag_mask_2),
    .io_from_addr_bits_tag_mask_3(Coalscer_io_from_addr_bits_tag_mask_3),
    .io_from_addr_bits_tag_mask_4(Coalscer_io_from_addr_bits_tag_mask_4),
    .io_from_addr_bits_tag_mask_5(Coalscer_io_from_addr_bits_tag_mask_5),
    .io_from_addr_bits_tag_mask_6(Coalscer_io_from_addr_bits_tag_mask_6),
    .io_from_addr_bits_tag_mask_7(Coalscer_io_from_addr_bits_tag_mask_7),
    .io_from_addr_bits_tag_unsigned(Coalscer_io_from_addr_bits_tag_unsigned),
    .io_from_addr_bits_tag_isvec(Coalscer_io_from_addr_bits_tag_isvec),
    .io_from_addr_bits_tag_isWrite(Coalscer_io_from_addr_bits_tag_isWrite),
    .io_idx_entry(Coalscer_io_idx_entry),
    .io_from_dcache_ready(Coalscer_io_from_dcache_ready),
    .io_from_dcache_valid(Coalscer_io_from_dcache_valid),
    .io_from_dcache_bits_instrId(Coalscer_io_from_dcache_bits_instrId),
    .io_from_dcache_bits_data_0(Coalscer_io_from_dcache_bits_data_0),
    .io_from_dcache_bits_data_1(Coalscer_io_from_dcache_bits_data_1),
    .io_from_dcache_bits_data_2(Coalscer_io_from_dcache_bits_data_2),
    .io_from_dcache_bits_data_3(Coalscer_io_from_dcache_bits_data_3),
    .io_from_dcache_bits_data_4(Coalscer_io_from_dcache_bits_data_4),
    .io_from_dcache_bits_data_5(Coalscer_io_from_dcache_bits_data_5),
    .io_from_dcache_bits_data_6(Coalscer_io_from_dcache_bits_data_6),
    .io_from_dcache_bits_data_7(Coalscer_io_from_dcache_bits_data_7),
    .io_from_dcache_bits_activeMask_0(Coalscer_io_from_dcache_bits_activeMask_0),
    .io_from_dcache_bits_activeMask_1(Coalscer_io_from_dcache_bits_activeMask_1),
    .io_from_dcache_bits_activeMask_2(Coalscer_io_from_dcache_bits_activeMask_2),
    .io_from_dcache_bits_activeMask_3(Coalscer_io_from_dcache_bits_activeMask_3),
    .io_from_dcache_bits_activeMask_4(Coalscer_io_from_dcache_bits_activeMask_4),
    .io_from_dcache_bits_activeMask_5(Coalscer_io_from_dcache_bits_activeMask_5),
    .io_from_dcache_bits_activeMask_6(Coalscer_io_from_dcache_bits_activeMask_6),
    .io_from_dcache_bits_activeMask_7(Coalscer_io_from_dcache_bits_activeMask_7),
    .io_to_pipe_ready(Coalscer_io_to_pipe_ready),
    .io_to_pipe_valid(Coalscer_io_to_pipe_valid),
    .io_to_pipe_bits_tag_warp_id(Coalscer_io_to_pipe_bits_tag_warp_id),
    .io_to_pipe_bits_tag_wfd(Coalscer_io_to_pipe_bits_tag_wfd),
    .io_to_pipe_bits_tag_wxd(Coalscer_io_to_pipe_bits_tag_wxd),
    .io_to_pipe_bits_tag_reg_idxw(Coalscer_io_to_pipe_bits_tag_reg_idxw),
    .io_to_pipe_bits_tag_mask_0(Coalscer_io_to_pipe_bits_tag_mask_0),
    .io_to_pipe_bits_tag_mask_1(Coalscer_io_to_pipe_bits_tag_mask_1),
    .io_to_pipe_bits_tag_mask_2(Coalscer_io_to_pipe_bits_tag_mask_2),
    .io_to_pipe_bits_tag_mask_3(Coalscer_io_to_pipe_bits_tag_mask_3),
    .io_to_pipe_bits_tag_mask_4(Coalscer_io_to_pipe_bits_tag_mask_4),
    .io_to_pipe_bits_tag_mask_5(Coalscer_io_to_pipe_bits_tag_mask_5),
    .io_to_pipe_bits_tag_mask_6(Coalscer_io_to_pipe_bits_tag_mask_6),
    .io_to_pipe_bits_tag_mask_7(Coalscer_io_to_pipe_bits_tag_mask_7),
    .io_to_pipe_bits_tag_isWrite(Coalscer_io_to_pipe_bits_tag_isWrite),
    .io_to_pipe_bits_data_0(Coalscer_io_to_pipe_bits_data_0),
    .io_to_pipe_bits_data_1(Coalscer_io_to_pipe_bits_data_1),
    .io_to_pipe_bits_data_2(Coalscer_io_to_pipe_bits_data_2),
    .io_to_pipe_bits_data_3(Coalscer_io_to_pipe_bits_data_3),
    .io_to_pipe_bits_data_4(Coalscer_io_to_pipe_bits_data_4),
    .io_to_pipe_bits_data_5(Coalscer_io_to_pipe_bits_data_5),
    .io_to_pipe_bits_data_6(Coalscer_io_to_pipe_bits_data_6),
    .io_to_pipe_bits_data_7(Coalscer_io_to_pipe_bits_data_7)
  );
  ShiftBoard ShiftBoard ( // @[LSU.scala 356:51]
    .clock(ShiftBoard_clock),
    .reset(ShiftBoard_reset),
    .io_left(ShiftBoard_io_left),
    .io_right(ShiftBoard_io_right),
    .io_full(ShiftBoard_io_full),
    .io_empty(ShiftBoard_io_empty)
  );
  ShiftBoard ShiftBoard_1 ( // @[LSU.scala 356:51]
    .clock(ShiftBoard_1_clock),
    .reset(ShiftBoard_1_reset),
    .io_left(ShiftBoard_1_io_left),
    .io_right(ShiftBoard_1_io_right),
    .io_full(ShiftBoard_1_io_full),
    .io_empty(ShiftBoard_1_io_empty)
  );
  ShiftBoard ShiftBoard_2 ( // @[LSU.scala 356:51]
    .clock(ShiftBoard_2_clock),
    .reset(ShiftBoard_2_reset),
    .io_left(ShiftBoard_2_io_left),
    .io_right(ShiftBoard_2_io_right),
    .io_full(ShiftBoard_2_io_full),
    .io_empty(ShiftBoard_2_io_empty)
  );
  ShiftBoard ShiftBoard_3 ( // @[LSU.scala 356:51]
    .clock(ShiftBoard_3_clock),
    .reset(ShiftBoard_3_reset),
    .io_left(ShiftBoard_3_io_left),
    .io_right(ShiftBoard_3_io_right),
    .io_full(ShiftBoard_3_io_full),
    .io_empty(ShiftBoard_3_io_empty)
  );
  assign io_lsu_req_ready = _GEN_3 ? 1'h0 : InputFIFO_io_enq_ready; // @[LSU.scala 362:24]
  assign io_dcache_rsp_ready = rspArbiter_io_in_0_ready; // @[LSU.scala 346:23]
  assign io_lsu_rsp_valid = Coalscer_io_to_pipe_valid; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_warp_id = Coalscer_io_to_pipe_bits_tag_warp_id; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_wfd = Coalscer_io_to_pipe_bits_tag_wfd; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_wxd = Coalscer_io_to_pipe_bits_tag_wxd; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_reg_idxw = Coalscer_io_to_pipe_bits_tag_reg_idxw; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_0 = Coalscer_io_to_pipe_bits_tag_mask_0; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_1 = Coalscer_io_to_pipe_bits_tag_mask_1; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_2 = Coalscer_io_to_pipe_bits_tag_mask_2; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_3 = Coalscer_io_to_pipe_bits_tag_mask_3; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_4 = Coalscer_io_to_pipe_bits_tag_mask_4; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_5 = Coalscer_io_to_pipe_bits_tag_mask_5; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_6 = Coalscer_io_to_pipe_bits_tag_mask_6; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_mask_7 = Coalscer_io_to_pipe_bits_tag_mask_7; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_tag_isWrite = Coalscer_io_to_pipe_bits_tag_isWrite; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_0 = Coalscer_io_to_pipe_bits_data_0; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_1 = Coalscer_io_to_pipe_bits_data_1; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_2 = Coalscer_io_to_pipe_bits_data_2; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_3 = Coalscer_io_to_pipe_bits_data_3; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_4 = Coalscer_io_to_pipe_bits_data_4; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_5 = Coalscer_io_to_pipe_bits_data_5; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_6 = Coalscer_io_to_pipe_bits_data_6; // @[LSU.scala 354:14]
  assign io_lsu_rsp_bits_data_7 = Coalscer_io_to_pipe_bits_data_7; // @[LSU.scala 354:14]
  assign io_dcache_req_valid = AddrCalc_io_to_dcache_valid; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_instrId = AddrCalc_io_to_dcache_bits_instrId; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_isWrite = AddrCalc_io_to_dcache_bits_isWrite; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_tag = AddrCalc_io_to_dcache_bits_tag; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_setIdx = AddrCalc_io_to_dcache_bits_setIdx; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_0_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_0_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_0_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_0_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_1_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_1_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_1_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_1_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_2_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_2_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_2_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_2_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_3_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_3_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_3_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_3_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_4_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_4_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_4_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_4_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_5_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_5_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_5_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_5_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_6_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_6_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_6_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_6_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_7_activeMask = AddrCalc_io_to_dcache_bits_perLaneAddr_7_activeMask; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_perLaneAddr_7_blockOffset = AddrCalc_io_to_dcache_bits_perLaneAddr_7_blockOffset; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_0 = AddrCalc_io_to_dcache_bits_data_0; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_1 = AddrCalc_io_to_dcache_bits_data_1; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_2 = AddrCalc_io_to_dcache_bits_data_2; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_3 = AddrCalc_io_to_dcache_bits_data_3; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_4 = AddrCalc_io_to_dcache_bits_data_4; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_5 = AddrCalc_io_to_dcache_bits_data_5; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_6 = AddrCalc_io_to_dcache_bits_data_6; // @[LSU.scala 341:17]
  assign io_dcache_req_bits_data_7 = AddrCalc_io_to_dcache_bits_data_7; // @[LSU.scala 341:17]
  assign io_shared_req_valid = AddrCalc_io_to_shared_valid; // @[LSU.scala 342:17]
  assign io_shared_req_bits_instrId = AddrCalc_io_to_shared_bits_instrId; // @[LSU.scala 342:17]
  assign io_shared_req_bits_isWrite = AddrCalc_io_to_shared_bits_isWrite; // @[LSU.scala 342:17]
  assign io_shared_req_bits_setIdx = AddrCalc_io_to_shared_bits_setIdx; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_0_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_0_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_0_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_0_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_1_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_1_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_1_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_1_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_2_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_2_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_2_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_2_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_3_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_3_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_3_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_3_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_4_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_4_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_4_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_4_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_5_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_5_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_5_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_5_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_6_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_6_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_6_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_6_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_7_activeMask = AddrCalc_io_to_shared_bits_perLaneAddr_7_activeMask; // @[LSU.scala 342:17]
  assign io_shared_req_bits_perLaneAddr_7_blockOffset = AddrCalc_io_to_shared_bits_perLaneAddr_7_blockOffset; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_0 = AddrCalc_io_to_shared_bits_data_0; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_1 = AddrCalc_io_to_shared_bits_data_1; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_2 = AddrCalc_io_to_shared_bits_data_2; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_3 = AddrCalc_io_to_shared_bits_data_3; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_4 = AddrCalc_io_to_shared_bits_data_4; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_5 = AddrCalc_io_to_shared_bits_data_5; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_6 = AddrCalc_io_to_shared_bits_data_6; // @[LSU.scala 342:17]
  assign io_shared_req_bits_data_7 = AddrCalc_io_to_shared_bits_data_7; // @[LSU.scala 342:17]
  assign io_shared_rsp_ready = rspArbiter_io_in_1_ready; // @[LSU.scala 345:23]
  assign io_fence_end = {io_fence_end_hi,io_fence_end_lo}; // @[LSU.scala 361:59]
  assign InputFIFO_clock = clock;
  assign InputFIFO_reset = reset;
  assign InputFIFO_io_enq_valid = _GEN_3 ? 1'h0 : io_lsu_req_valid; // @[LSU.scala 363:30]
  assign InputFIFO_io_enq_bits_in1_0 = io_lsu_req_bits_in1_0; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_1 = io_lsu_req_bits_in1_1; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_2 = io_lsu_req_bits_in1_2; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_3 = io_lsu_req_bits_in1_3; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_4 = io_lsu_req_bits_in1_4; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_5 = io_lsu_req_bits_in1_5; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_6 = io_lsu_req_bits_in1_6; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in1_7 = io_lsu_req_bits_in1_7; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_0 = io_lsu_req_bits_in2_0; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_1 = io_lsu_req_bits_in2_1; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_2 = io_lsu_req_bits_in2_2; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_3 = io_lsu_req_bits_in2_3; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_4 = io_lsu_req_bits_in2_4; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_5 = io_lsu_req_bits_in2_5; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_6 = io_lsu_req_bits_in2_6; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in2_7 = io_lsu_req_bits_in2_7; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_0 = io_lsu_req_bits_in3_0; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_1 = io_lsu_req_bits_in3_1; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_2 = io_lsu_req_bits_in3_2; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_3 = io_lsu_req_bits_in3_3; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_4 = io_lsu_req_bits_in3_4; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_5 = io_lsu_req_bits_in3_5; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_6 = io_lsu_req_bits_in3_6; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_in3_7 = io_lsu_req_bits_in3_7; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_0 = io_lsu_req_bits_mask_0; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_1 = io_lsu_req_bits_mask_1; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_2 = io_lsu_req_bits_mask_2; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_3 = io_lsu_req_bits_mask_3; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_4 = io_lsu_req_bits_mask_4; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_5 = io_lsu_req_bits_mask_5; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_6 = io_lsu_req_bits_mask_6; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_mask_7 = io_lsu_req_bits_mask_7; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_inst = io_lsu_req_bits_ctrl_inst; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_wid = io_lsu_req_bits_ctrl_wid; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_fp = io_lsu_req_bits_ctrl_fp; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_branch = io_lsu_req_bits_ctrl_branch; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_simt_stack = io_lsu_req_bits_ctrl_simt_stack; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_simt_stack_op = io_lsu_req_bits_ctrl_simt_stack_op; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_barrier = io_lsu_req_bits_ctrl_barrier; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_csr = io_lsu_req_bits_ctrl_csr; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_reverse = io_lsu_req_bits_ctrl_reverse; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_isvec = io_lsu_req_bits_ctrl_isvec; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_mem_unsigned = io_lsu_req_bits_ctrl_mem_unsigned; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_alu_fn = io_lsu_req_bits_ctrl_alu_fn; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_mem = io_lsu_req_bits_ctrl_mem; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_mem_cmd = io_lsu_req_bits_ctrl_mem_cmd; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_mop = io_lsu_req_bits_ctrl_mop; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_reg_idxw = io_lsu_req_bits_ctrl_reg_idxw; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_wfd = io_lsu_req_bits_ctrl_wfd; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_fence = io_lsu_req_bits_ctrl_fence; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_sfu = io_lsu_req_bits_ctrl_sfu; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_readmask = io_lsu_req_bits_ctrl_readmask; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_writemask = io_lsu_req_bits_ctrl_writemask; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_wxd = io_lsu_req_bits_ctrl_wxd; // @[LSU.scala 337:20]
  assign InputFIFO_io_enq_bits_ctrl_pc = io_lsu_req_bits_ctrl_pc; // @[LSU.scala 337:20]
  assign InputFIFO_io_deq_ready = AddrCalc_io_from_fifo_ready; // @[LSU.scala 340:25]
  assign AddrCalc_clock = clock;
  assign AddrCalc_reset = reset;
  assign AddrCalc_io_from_fifo_valid = InputFIFO_io_deq_valid; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_0 = InputFIFO_io_deq_bits_in1_0; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_1 = InputFIFO_io_deq_bits_in1_1; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_2 = InputFIFO_io_deq_bits_in1_2; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_3 = InputFIFO_io_deq_bits_in1_3; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_4 = InputFIFO_io_deq_bits_in1_4; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_5 = InputFIFO_io_deq_bits_in1_5; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_6 = InputFIFO_io_deq_bits_in1_6; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in1_7 = InputFIFO_io_deq_bits_in1_7; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_0 = InputFIFO_io_deq_bits_in2_0; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_1 = InputFIFO_io_deq_bits_in2_1; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_2 = InputFIFO_io_deq_bits_in2_2; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_3 = InputFIFO_io_deq_bits_in2_3; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_4 = InputFIFO_io_deq_bits_in2_4; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_5 = InputFIFO_io_deq_bits_in2_5; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_6 = InputFIFO_io_deq_bits_in2_6; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in2_7 = InputFIFO_io_deq_bits_in2_7; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_0 = InputFIFO_io_deq_bits_in3_0; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_1 = InputFIFO_io_deq_bits_in3_1; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_2 = InputFIFO_io_deq_bits_in3_2; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_3 = InputFIFO_io_deq_bits_in3_3; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_4 = InputFIFO_io_deq_bits_in3_4; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_5 = InputFIFO_io_deq_bits_in3_5; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_6 = InputFIFO_io_deq_bits_in3_6; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_in3_7 = InputFIFO_io_deq_bits_in3_7; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_0 = InputFIFO_io_deq_bits_mask_0; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_1 = InputFIFO_io_deq_bits_mask_1; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_2 = InputFIFO_io_deq_bits_mask_2; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_3 = InputFIFO_io_deq_bits_mask_3; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_4 = InputFIFO_io_deq_bits_mask_4; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_5 = InputFIFO_io_deq_bits_mask_5; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_6 = InputFIFO_io_deq_bits_mask_6; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_mask_7 = InputFIFO_io_deq_bits_mask_7; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_wid = InputFIFO_io_deq_bits_ctrl_wid; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_isvec = InputFIFO_io_deq_bits_ctrl_isvec; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_mem_unsigned = InputFIFO_io_deq_bits_ctrl_mem_unsigned; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_mem_cmd = InputFIFO_io_deq_bits_ctrl_mem_cmd; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_mop = InputFIFO_io_deq_bits_ctrl_mop; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_reg_idxw = InputFIFO_io_deq_bits_ctrl_reg_idxw; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_wfd = InputFIFO_io_deq_bits_ctrl_wfd; // @[LSU.scala 340:25]
  assign AddrCalc_io_from_fifo_bits_ctrl_wxd = InputFIFO_io_deq_bits_ctrl_wxd; // @[LSU.scala 340:25]
  assign AddrCalc_io_to_mshr_ready = Coalscer_io_from_addr_ready; // @[LSU.scala 352:25]
  assign AddrCalc_io_idx_entry = Coalscer_io_idx_entry; // @[LSU.scala 353:24]
  assign AddrCalc_io_to_dcache_ready = io_dcache_req_ready; // @[LSU.scala 341:17]
  assign AddrCalc_io_to_shared_ready = io_shared_req_ready; // @[LSU.scala 342:17]
  assign rspArbiter_io_in_0_valid = io_dcache_rsp_valid; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_instrId = io_dcache_rsp_bits_instrId; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_0 = io_dcache_rsp_bits_data_0; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_1 = io_dcache_rsp_bits_data_1; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_2 = io_dcache_rsp_bits_data_2; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_3 = io_dcache_rsp_bits_data_3; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_4 = io_dcache_rsp_bits_data_4; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_5 = io_dcache_rsp_bits_data_5; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_6 = io_dcache_rsp_bits_data_6; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_data_7 = io_dcache_rsp_bits_data_7; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_0 = io_dcache_rsp_bits_activeMask_0; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_1 = io_dcache_rsp_bits_activeMask_1; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_2 = io_dcache_rsp_bits_activeMask_2; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_3 = io_dcache_rsp_bits_activeMask_3; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_4 = io_dcache_rsp_bits_activeMask_4; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_5 = io_dcache_rsp_bits_activeMask_5; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_6 = io_dcache_rsp_bits_activeMask_6; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_0_bits_activeMask_7 = io_dcache_rsp_bits_activeMask_7; // @[LSU.scala 346:23]
  assign rspArbiter_io_in_1_valid = io_shared_rsp_valid; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_instrId = io_shared_rsp_bits_instrId; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_0 = io_shared_rsp_bits_data_0; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_1 = io_shared_rsp_bits_data_1; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_2 = io_shared_rsp_bits_data_2; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_3 = io_shared_rsp_bits_data_3; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_4 = io_shared_rsp_bits_data_4; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_5 = io_shared_rsp_bits_data_5; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_6 = io_shared_rsp_bits_data_6; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_data_7 = io_shared_rsp_bits_data_7; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_0 = io_shared_rsp_bits_activeMask_0; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_1 = io_shared_rsp_bits_activeMask_1; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_2 = io_shared_rsp_bits_activeMask_2; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_3 = io_shared_rsp_bits_activeMask_3; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_4 = io_shared_rsp_bits_activeMask_4; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_5 = io_shared_rsp_bits_activeMask_5; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_6 = io_shared_rsp_bits_activeMask_6; // @[LSU.scala 345:23]
  assign rspArbiter_io_in_1_bits_activeMask_7 = io_shared_rsp_bits_activeMask_7; // @[LSU.scala 345:23]
  assign rspArbiter_io_out_ready = Coalscer_io_from_dcache_ready; // @[LSU.scala 351:27]
  assign Coalscer_clock = clock;
  assign Coalscer_reset = reset;
  assign Coalscer_io_from_addr_valid = AddrCalc_io_to_mshr_valid; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_warp_id = AddrCalc_io_to_mshr_bits_tag_warp_id; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_wfd = AddrCalc_io_to_mshr_bits_tag_wfd; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_wxd = AddrCalc_io_to_mshr_bits_tag_wxd; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_reg_idxw = AddrCalc_io_to_mshr_bits_tag_reg_idxw; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_0 = AddrCalc_io_to_mshr_bits_tag_mask_0; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_1 = AddrCalc_io_to_mshr_bits_tag_mask_1; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_2 = AddrCalc_io_to_mshr_bits_tag_mask_2; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_3 = AddrCalc_io_to_mshr_bits_tag_mask_3; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_4 = AddrCalc_io_to_mshr_bits_tag_mask_4; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_5 = AddrCalc_io_to_mshr_bits_tag_mask_5; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_6 = AddrCalc_io_to_mshr_bits_tag_mask_6; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_mask_7 = AddrCalc_io_to_mshr_bits_tag_mask_7; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_unsigned = AddrCalc_io_to_mshr_bits_tag_unsigned; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_isvec = AddrCalc_io_to_mshr_bits_tag_isvec; // @[LSU.scala 352:25]
  assign Coalscer_io_from_addr_bits_tag_isWrite = AddrCalc_io_to_mshr_bits_tag_isWrite; // @[LSU.scala 352:25]
  assign Coalscer_io_from_dcache_valid = rspArbiter_io_out_valid; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_instrId = rspArbiter_io_out_bits_instrId; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_0 = rspArbiter_io_out_bits_data_0; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_1 = rspArbiter_io_out_bits_data_1; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_2 = rspArbiter_io_out_bits_data_2; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_3 = rspArbiter_io_out_bits_data_3; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_4 = rspArbiter_io_out_bits_data_4; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_5 = rspArbiter_io_out_bits_data_5; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_6 = rspArbiter_io_out_bits_data_6; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_data_7 = rspArbiter_io_out_bits_data_7; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_0 = rspArbiter_io_out_bits_activeMask_0; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_1 = rspArbiter_io_out_bits_activeMask_1; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_2 = rspArbiter_io_out_bits_activeMask_2; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_3 = rspArbiter_io_out_bits_activeMask_3; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_4 = rspArbiter_io_out_bits_activeMask_4; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_5 = rspArbiter_io_out_bits_activeMask_5; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_6 = rspArbiter_io_out_bits_activeMask_6; // @[LSU.scala 351:27]
  assign Coalscer_io_from_dcache_bits_activeMask_7 = rspArbiter_io_out_bits_activeMask_7; // @[LSU.scala 351:27]
  assign Coalscer_io_to_pipe_ready = io_lsu_rsp_ready; // @[LSU.scala 354:14]
  assign ShiftBoard_clock = clock;
  assign ShiftBoard_reset = reset;
  assign ShiftBoard_io_left = _shiftBoard_0_left_T & io_lsu_req_bits_ctrl_wid == 2'h0; // @[LSU.scala 358:29]
  assign ShiftBoard_io_right = _shiftBoard_0_right_T & io_lsu_rsp_bits_tag_warp_id == 2'h0; // @[LSU.scala 359:30]
  assign ShiftBoard_1_clock = clock;
  assign ShiftBoard_1_reset = reset;
  assign ShiftBoard_1_io_left = _shiftBoard_0_left_T & io_lsu_req_bits_ctrl_wid == 2'h1; // @[LSU.scala 358:29]
  assign ShiftBoard_1_io_right = _shiftBoard_0_right_T & io_lsu_rsp_bits_tag_warp_id == 2'h1; // @[LSU.scala 359:30]
  assign ShiftBoard_2_clock = clock;
  assign ShiftBoard_2_reset = reset;
  assign ShiftBoard_2_io_left = _shiftBoard_0_left_T & io_lsu_req_bits_ctrl_wid == 2'h2; // @[LSU.scala 358:29]
  assign ShiftBoard_2_io_right = _shiftBoard_0_right_T & io_lsu_rsp_bits_tag_warp_id == 2'h2; // @[LSU.scala 359:30]
  assign ShiftBoard_3_clock = clock;
  assign ShiftBoard_3_reset = reset;
  assign ShiftBoard_3_io_left = _shiftBoard_0_left_T & io_lsu_req_bits_ctrl_wid == 2'h3; // @[LSU.scala 358:29]
  assign ShiftBoard_3_io_right = _shiftBoard_0_right_T & io_lsu_rsp_bits_tag_warp_id == 2'h3; // @[LSU.scala 359:30]
endmodule
module Queue_44(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_in1_0,
  input  [31:0] io_enq_bits_in1_1,
  input  [31:0] io_enq_bits_in1_2,
  input  [31:0] io_enq_bits_in1_3,
  input  [31:0] io_enq_bits_in1_4,
  input  [31:0] io_enq_bits_in1_5,
  input  [31:0] io_enq_bits_in1_6,
  input  [31:0] io_enq_bits_in1_7,
  input  [31:0] io_enq_bits_in2_0,
  input  [31:0] io_enq_bits_in2_1,
  input  [31:0] io_enq_bits_in2_2,
  input  [31:0] io_enq_bits_in2_3,
  input  [31:0] io_enq_bits_in2_4,
  input  [31:0] io_enq_bits_in2_5,
  input  [31:0] io_enq_bits_in2_6,
  input  [31:0] io_enq_bits_in2_7,
  input         io_enq_bits_mask_0,
  input         io_enq_bits_mask_1,
  input         io_enq_bits_mask_2,
  input         io_enq_bits_mask_3,
  input         io_enq_bits_mask_4,
  input         io_enq_bits_mask_5,
  input         io_enq_bits_mask_6,
  input         io_enq_bits_mask_7,
  input  [1:0]  io_enq_bits_ctrl_wid,
  input         io_enq_bits_ctrl_fp,
  input         io_enq_bits_ctrl_reverse,
  input         io_enq_bits_ctrl_isvec,
  input  [5:0]  io_enq_bits_ctrl_alu_fn,
  input  [4:0]  io_enq_bits_ctrl_reg_idxw,
  input         io_enq_bits_ctrl_wfd,
  input         io_enq_bits_ctrl_wxd,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_in1_0,
  output [31:0] io_deq_bits_in1_1,
  output [31:0] io_deq_bits_in1_2,
  output [31:0] io_deq_bits_in1_3,
  output [31:0] io_deq_bits_in1_4,
  output [31:0] io_deq_bits_in1_5,
  output [31:0] io_deq_bits_in1_6,
  output [31:0] io_deq_bits_in1_7,
  output [31:0] io_deq_bits_in2_0,
  output [31:0] io_deq_bits_in2_1,
  output [31:0] io_deq_bits_in2_2,
  output [31:0] io_deq_bits_in2_3,
  output [31:0] io_deq_bits_in2_4,
  output [31:0] io_deq_bits_in2_5,
  output [31:0] io_deq_bits_in2_6,
  output [31:0] io_deq_bits_in2_7,
  output        io_deq_bits_mask_0,
  output        io_deq_bits_mask_1,
  output        io_deq_bits_mask_2,
  output        io_deq_bits_mask_3,
  output        io_deq_bits_mask_4,
  output        io_deq_bits_mask_5,
  output        io_deq_bits_mask_6,
  output        io_deq_bits_mask_7,
  output [1:0]  io_deq_bits_ctrl_wid,
  output        io_deq_bits_ctrl_fp,
  output        io_deq_bits_ctrl_reverse,
  output        io_deq_bits_ctrl_isvec,
  output [5:0]  io_deq_bits_ctrl_alu_fn,
  output [4:0]  io_deq_bits_ctrl_reg_idxw,
  output        io_deq_bits_ctrl_wfd,
  output        io_deq_bits_ctrl_wxd
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_in1_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in1_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in1_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in1_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_in2_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_in2_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_in2_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_mask_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_ctrl_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_fp [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_fp_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_reverse [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reverse_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_isvec [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_isvec_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] ram_ctrl_alu_fn [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [5:0] ram_ctrl_alu_fn_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_ctrl_alu_fn_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_alu_fn_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_ctrl_reg_idxw [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_reg_idxw_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wfd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wfd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_ctrl_wxd [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_ctrl_wxd_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_in1_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_0_io_deq_bits_MPORT_data = ram_in1_0[ram_in1_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_0_MPORT_data = io_enq_bits_in1_0;
  assign ram_in1_0_MPORT_addr = 1'h0;
  assign ram_in1_0_MPORT_mask = 1'h1;
  assign ram_in1_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_1_io_deq_bits_MPORT_data = ram_in1_1[ram_in1_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_1_MPORT_data = io_enq_bits_in1_1;
  assign ram_in1_1_MPORT_addr = 1'h0;
  assign ram_in1_1_MPORT_mask = 1'h1;
  assign ram_in1_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_2_io_deq_bits_MPORT_data = ram_in1_2[ram_in1_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_2_MPORT_data = io_enq_bits_in1_2;
  assign ram_in1_2_MPORT_addr = 1'h0;
  assign ram_in1_2_MPORT_mask = 1'h1;
  assign ram_in1_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_3_io_deq_bits_MPORT_data = ram_in1_3[ram_in1_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_3_MPORT_data = io_enq_bits_in1_3;
  assign ram_in1_3_MPORT_addr = 1'h0;
  assign ram_in1_3_MPORT_mask = 1'h1;
  assign ram_in1_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_4_io_deq_bits_MPORT_data = ram_in1_4[ram_in1_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_4_MPORT_data = io_enq_bits_in1_4;
  assign ram_in1_4_MPORT_addr = 1'h0;
  assign ram_in1_4_MPORT_mask = 1'h1;
  assign ram_in1_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_5_io_deq_bits_MPORT_data = ram_in1_5[ram_in1_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_5_MPORT_data = io_enq_bits_in1_5;
  assign ram_in1_5_MPORT_addr = 1'h0;
  assign ram_in1_5_MPORT_mask = 1'h1;
  assign ram_in1_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_6_io_deq_bits_MPORT_data = ram_in1_6[ram_in1_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_6_MPORT_data = io_enq_bits_in1_6;
  assign ram_in1_6_MPORT_addr = 1'h0;
  assign ram_in1_6_MPORT_mask = 1'h1;
  assign ram_in1_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in1_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in1_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in1_7_io_deq_bits_MPORT_data = ram_in1_7[ram_in1_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in1_7_MPORT_data = io_enq_bits_in1_7;
  assign ram_in1_7_MPORT_addr = 1'h0;
  assign ram_in1_7_MPORT_mask = 1'h1;
  assign ram_in1_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_0_io_deq_bits_MPORT_data = ram_in2_0[ram_in2_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_0_MPORT_data = io_enq_bits_in2_0;
  assign ram_in2_0_MPORT_addr = 1'h0;
  assign ram_in2_0_MPORT_mask = 1'h1;
  assign ram_in2_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_1_io_deq_bits_MPORT_data = ram_in2_1[ram_in2_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_1_MPORT_data = io_enq_bits_in2_1;
  assign ram_in2_1_MPORT_addr = 1'h0;
  assign ram_in2_1_MPORT_mask = 1'h1;
  assign ram_in2_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_2_io_deq_bits_MPORT_data = ram_in2_2[ram_in2_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_2_MPORT_data = io_enq_bits_in2_2;
  assign ram_in2_2_MPORT_addr = 1'h0;
  assign ram_in2_2_MPORT_mask = 1'h1;
  assign ram_in2_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_3_io_deq_bits_MPORT_data = ram_in2_3[ram_in2_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_3_MPORT_data = io_enq_bits_in2_3;
  assign ram_in2_3_MPORT_addr = 1'h0;
  assign ram_in2_3_MPORT_mask = 1'h1;
  assign ram_in2_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_4_io_deq_bits_MPORT_data = ram_in2_4[ram_in2_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_4_MPORT_data = io_enq_bits_in2_4;
  assign ram_in2_4_MPORT_addr = 1'h0;
  assign ram_in2_4_MPORT_mask = 1'h1;
  assign ram_in2_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_5_io_deq_bits_MPORT_data = ram_in2_5[ram_in2_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_5_MPORT_data = io_enq_bits_in2_5;
  assign ram_in2_5_MPORT_addr = 1'h0;
  assign ram_in2_5_MPORT_mask = 1'h1;
  assign ram_in2_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_6_io_deq_bits_MPORT_data = ram_in2_6[ram_in2_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_6_MPORT_data = io_enq_bits_in2_6;
  assign ram_in2_6_MPORT_addr = 1'h0;
  assign ram_in2_6_MPORT_mask = 1'h1;
  assign ram_in2_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_in2_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_in2_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_in2_7_io_deq_bits_MPORT_data = ram_in2_7[ram_in2_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_in2_7_MPORT_data = io_enq_bits_in2_7;
  assign ram_in2_7_MPORT_addr = 1'h0;
  assign ram_in2_7_MPORT_mask = 1'h1;
  assign ram_in2_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_0_io_deq_bits_MPORT_data = ram_mask_0[ram_mask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_0_MPORT_data = io_enq_bits_mask_0;
  assign ram_mask_0_MPORT_addr = 1'h0;
  assign ram_mask_0_MPORT_mask = 1'h1;
  assign ram_mask_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_1_io_deq_bits_MPORT_data = ram_mask_1[ram_mask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_1_MPORT_data = io_enq_bits_mask_1;
  assign ram_mask_1_MPORT_addr = 1'h0;
  assign ram_mask_1_MPORT_mask = 1'h1;
  assign ram_mask_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_2_io_deq_bits_MPORT_data = ram_mask_2[ram_mask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_2_MPORT_data = io_enq_bits_mask_2;
  assign ram_mask_2_MPORT_addr = 1'h0;
  assign ram_mask_2_MPORT_mask = 1'h1;
  assign ram_mask_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_3_io_deq_bits_MPORT_data = ram_mask_3[ram_mask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_3_MPORT_data = io_enq_bits_mask_3;
  assign ram_mask_3_MPORT_addr = 1'h0;
  assign ram_mask_3_MPORT_mask = 1'h1;
  assign ram_mask_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_4_io_deq_bits_MPORT_data = ram_mask_4[ram_mask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_4_MPORT_data = io_enq_bits_mask_4;
  assign ram_mask_4_MPORT_addr = 1'h0;
  assign ram_mask_4_MPORT_mask = 1'h1;
  assign ram_mask_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_5_io_deq_bits_MPORT_data = ram_mask_5[ram_mask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_5_MPORT_data = io_enq_bits_mask_5;
  assign ram_mask_5_MPORT_addr = 1'h0;
  assign ram_mask_5_MPORT_mask = 1'h1;
  assign ram_mask_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_6_io_deq_bits_MPORT_data = ram_mask_6[ram_mask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_6_MPORT_data = io_enq_bits_mask_6;
  assign ram_mask_6_MPORT_addr = 1'h0;
  assign ram_mask_6_MPORT_mask = 1'h1;
  assign ram_mask_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_7_io_deq_bits_MPORT_data = ram_mask_7[ram_mask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_7_MPORT_data = io_enq_bits_mask_7;
  assign ram_mask_7_MPORT_addr = 1'h0;
  assign ram_mask_7_MPORT_mask = 1'h1;
  assign ram_mask_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wid_io_deq_bits_MPORT_data = ram_ctrl_wid[ram_ctrl_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wid_MPORT_data = io_enq_bits_ctrl_wid;
  assign ram_ctrl_wid_MPORT_addr = 1'h0;
  assign ram_ctrl_wid_MPORT_mask = 1'h1;
  assign ram_ctrl_wid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_fp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_fp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_fp_io_deq_bits_MPORT_data = ram_ctrl_fp[ram_ctrl_fp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_fp_MPORT_data = io_enq_bits_ctrl_fp;
  assign ram_ctrl_fp_MPORT_addr = 1'h0;
  assign ram_ctrl_fp_MPORT_mask = 1'h1;
  assign ram_ctrl_fp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_reverse_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_reverse_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_reverse_io_deq_bits_MPORT_data = ram_ctrl_reverse[ram_ctrl_reverse_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_reverse_MPORT_data = io_enq_bits_ctrl_reverse;
  assign ram_ctrl_reverse_MPORT_addr = 1'h0;
  assign ram_ctrl_reverse_MPORT_mask = 1'h1;
  assign ram_ctrl_reverse_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_isvec_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_isvec_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_isvec_io_deq_bits_MPORT_data = ram_ctrl_isvec[ram_ctrl_isvec_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_isvec_MPORT_data = io_enq_bits_ctrl_isvec;
  assign ram_ctrl_isvec_MPORT_addr = 1'h0;
  assign ram_ctrl_isvec_MPORT_mask = 1'h1;
  assign ram_ctrl_isvec_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_alu_fn_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_alu_fn_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_alu_fn_io_deq_bits_MPORT_data = ram_ctrl_alu_fn[ram_ctrl_alu_fn_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_alu_fn_MPORT_data = io_enq_bits_ctrl_alu_fn;
  assign ram_ctrl_alu_fn_MPORT_addr = 1'h0;
  assign ram_ctrl_alu_fn_MPORT_mask = 1'h1;
  assign ram_ctrl_alu_fn_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_reg_idxw_io_deq_bits_MPORT_data = ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_reg_idxw_MPORT_data = io_enq_bits_ctrl_reg_idxw;
  assign ram_ctrl_reg_idxw_MPORT_addr = 1'h0;
  assign ram_ctrl_reg_idxw_MPORT_mask = 1'h1;
  assign ram_ctrl_reg_idxw_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wfd_io_deq_bits_MPORT_data = ram_ctrl_wfd[ram_ctrl_wfd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wfd_MPORT_data = io_enq_bits_ctrl_wfd;
  assign ram_ctrl_wfd_MPORT_addr = 1'h0;
  assign ram_ctrl_wfd_MPORT_mask = 1'h1;
  assign ram_ctrl_wfd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_ctrl_wxd_io_deq_bits_MPORT_data = ram_ctrl_wxd[ram_ctrl_wxd_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_ctrl_wxd_MPORT_data = io_enq_bits_ctrl_wxd;
  assign ram_ctrl_wxd_MPORT_addr = 1'h0;
  assign ram_ctrl_wxd_MPORT_mask = 1'h1;
  assign ram_ctrl_wxd_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_in1_0 = ram_in1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_1 = ram_in1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_2 = ram_in1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_3 = ram_in1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_4 = ram_in1_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_5 = ram_in1_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_6 = ram_in1_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in1_7 = ram_in1_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_0 = ram_in2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_1 = ram_in2_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_2 = ram_in2_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_3 = ram_in2_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_4 = ram_in2_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_5 = ram_in2_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_6 = ram_in2_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_in2_7 = ram_in2_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_0 = ram_mask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_1 = ram_mask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_2 = ram_mask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_3 = ram_mask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_4 = ram_mask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_5 = ram_mask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_6 = ram_mask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask_7 = ram_mask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_wid = ram_ctrl_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_fp = ram_ctrl_fp_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_reverse = ram_ctrl_reverse_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_isvec = ram_ctrl_isvec_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_alu_fn = ram_ctrl_alu_fn_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_reg_idxw = ram_ctrl_reg_idxw_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_wfd = ram_ctrl_wfd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_ctrl_wxd = ram_ctrl_wxd_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_in1_0_MPORT_en & ram_in1_0_MPORT_mask) begin
      ram_in1_0[ram_in1_0_MPORT_addr] <= ram_in1_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_1_MPORT_en & ram_in1_1_MPORT_mask) begin
      ram_in1_1[ram_in1_1_MPORT_addr] <= ram_in1_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_2_MPORT_en & ram_in1_2_MPORT_mask) begin
      ram_in1_2[ram_in1_2_MPORT_addr] <= ram_in1_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_3_MPORT_en & ram_in1_3_MPORT_mask) begin
      ram_in1_3[ram_in1_3_MPORT_addr] <= ram_in1_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_4_MPORT_en & ram_in1_4_MPORT_mask) begin
      ram_in1_4[ram_in1_4_MPORT_addr] <= ram_in1_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_5_MPORT_en & ram_in1_5_MPORT_mask) begin
      ram_in1_5[ram_in1_5_MPORT_addr] <= ram_in1_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_6_MPORT_en & ram_in1_6_MPORT_mask) begin
      ram_in1_6[ram_in1_6_MPORT_addr] <= ram_in1_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in1_7_MPORT_en & ram_in1_7_MPORT_mask) begin
      ram_in1_7[ram_in1_7_MPORT_addr] <= ram_in1_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_0_MPORT_en & ram_in2_0_MPORT_mask) begin
      ram_in2_0[ram_in2_0_MPORT_addr] <= ram_in2_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_1_MPORT_en & ram_in2_1_MPORT_mask) begin
      ram_in2_1[ram_in2_1_MPORT_addr] <= ram_in2_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_2_MPORT_en & ram_in2_2_MPORT_mask) begin
      ram_in2_2[ram_in2_2_MPORT_addr] <= ram_in2_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_3_MPORT_en & ram_in2_3_MPORT_mask) begin
      ram_in2_3[ram_in2_3_MPORT_addr] <= ram_in2_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_4_MPORT_en & ram_in2_4_MPORT_mask) begin
      ram_in2_4[ram_in2_4_MPORT_addr] <= ram_in2_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_5_MPORT_en & ram_in2_5_MPORT_mask) begin
      ram_in2_5[ram_in2_5_MPORT_addr] <= ram_in2_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_6_MPORT_en & ram_in2_6_MPORT_mask) begin
      ram_in2_6[ram_in2_6_MPORT_addr] <= ram_in2_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_in2_7_MPORT_en & ram_in2_7_MPORT_mask) begin
      ram_in2_7[ram_in2_7_MPORT_addr] <= ram_in2_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_0_MPORT_en & ram_mask_0_MPORT_mask) begin
      ram_mask_0[ram_mask_0_MPORT_addr] <= ram_mask_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_1_MPORT_en & ram_mask_1_MPORT_mask) begin
      ram_mask_1[ram_mask_1_MPORT_addr] <= ram_mask_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_2_MPORT_en & ram_mask_2_MPORT_mask) begin
      ram_mask_2[ram_mask_2_MPORT_addr] <= ram_mask_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_3_MPORT_en & ram_mask_3_MPORT_mask) begin
      ram_mask_3[ram_mask_3_MPORT_addr] <= ram_mask_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_4_MPORT_en & ram_mask_4_MPORT_mask) begin
      ram_mask_4[ram_mask_4_MPORT_addr] <= ram_mask_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_5_MPORT_en & ram_mask_5_MPORT_mask) begin
      ram_mask_5[ram_mask_5_MPORT_addr] <= ram_mask_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_6_MPORT_en & ram_mask_6_MPORT_mask) begin
      ram_mask_6[ram_mask_6_MPORT_addr] <= ram_mask_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_7_MPORT_en & ram_mask_7_MPORT_mask) begin
      ram_mask_7[ram_mask_7_MPORT_addr] <= ram_mask_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wid_MPORT_en & ram_ctrl_wid_MPORT_mask) begin
      ram_ctrl_wid[ram_ctrl_wid_MPORT_addr] <= ram_ctrl_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_fp_MPORT_en & ram_ctrl_fp_MPORT_mask) begin
      ram_ctrl_fp[ram_ctrl_fp_MPORT_addr] <= ram_ctrl_fp_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_reverse_MPORT_en & ram_ctrl_reverse_MPORT_mask) begin
      ram_ctrl_reverse[ram_ctrl_reverse_MPORT_addr] <= ram_ctrl_reverse_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_isvec_MPORT_en & ram_ctrl_isvec_MPORT_mask) begin
      ram_ctrl_isvec[ram_ctrl_isvec_MPORT_addr] <= ram_ctrl_isvec_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_alu_fn_MPORT_en & ram_ctrl_alu_fn_MPORT_mask) begin
      ram_ctrl_alu_fn[ram_ctrl_alu_fn_MPORT_addr] <= ram_ctrl_alu_fn_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_reg_idxw_MPORT_en & ram_ctrl_reg_idxw_MPORT_mask) begin
      ram_ctrl_reg_idxw[ram_ctrl_reg_idxw_MPORT_addr] <= ram_ctrl_reg_idxw_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wfd_MPORT_en & ram_ctrl_wfd_MPORT_mask) begin
      ram_ctrl_wfd[ram_ctrl_wfd_MPORT_addr] <= ram_ctrl_wfd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_ctrl_wxd_MPORT_en & ram_ctrl_wxd_MPORT_mask) begin
      ram_ctrl_wxd[ram_ctrl_wxd_MPORT_addr] <= ram_ctrl_wxd_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_0[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_1[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_2[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_3[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_4[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_5[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_6[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in1_7[initvar] = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_0[initvar] = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_1[initvar] = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_2[initvar] = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_3[initvar] = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_4[initvar] = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_5[initvar] = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_6[initvar] = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_in2_7[initvar] = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_0[initvar] = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_1[initvar] = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_2[initvar] = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_3[initvar] = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_4[initvar] = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_5[initvar] = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_6[initvar] = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_7[initvar] = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wid[initvar] = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_fp[initvar] = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_reverse[initvar] = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_isvec[initvar] = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_alu_fn[initvar] = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_reg_idxw[initvar] = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wfd[initvar] = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_ctrl_wxd[initvar] = _RAND_31[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  maybe_full = _RAND_32[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IntDivMod(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_a,
  input  [31:0] io_in_bits_d,
  input         io_in_bits_signed,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_q,
  output [31:0] io_out_bits_r
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[IntDivMod.scala 16:22]
  wire  aSign = io_in_bits_signed & io_in_bits_a[31]; // @[IntDivMod.scala 18:33]
  wire  dSign = io_in_bits_signed & io_in_bits_d[31]; // @[IntDivMod.scala 19:33]
  wire  _qSignReg_T = aSign ^ dSign; // @[IntDivMod.scala 20:34]
  wire  _qSignReg_T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  reg  qSignReg; // @[Reg.scala 16:16]
  reg  rSignReg; // @[Reg.scala 16:16]
  wire [31:0] _unsignedA_T = ~io_in_bits_a; // @[IntDivMod.scala 22:31]
  wire [31:0] _unsignedA_T_2 = _unsignedA_T + 32'h1; // @[IntDivMod.scala 22:54]
  wire [31:0] _unsignedD_T = ~io_in_bits_d; // @[IntDivMod.scala 23:31]
  wire [31:0] _unsignedD_T_2 = _unsignedD_T + 32'h1; // @[IntDivMod.scala 23:54]
  wire  overflow = aSign & ~(|io_in_bits_a[30:0]) & &io_in_bits_d; // @[IntDivMod.scala 25:100]
  wire  divByZero = io_in_bits_d == 32'h0; // @[IntDivMod.scala 26:32]
  reg [31:0] rawAReg; // @[Reg.scala 16:16]
  reg [31:0] unsignedAReg; // @[Reg.scala 16:16]
  reg [31:0] unsignedDReg; // @[Reg.scala 16:16]
  reg  overflowReg; // @[Reg.scala 16:16]
  reg  divByZeroReg; // @[Reg.scala 16:16]
  wire [4:0] _aLez_T_32 = unsignedAReg[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_33 = unsignedAReg[2] ? 5'h1d : _aLez_T_32; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_34 = unsignedAReg[3] ? 5'h1c : _aLez_T_33; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_35 = unsignedAReg[4] ? 5'h1b : _aLez_T_34; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_36 = unsignedAReg[5] ? 5'h1a : _aLez_T_35; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_37 = unsignedAReg[6] ? 5'h19 : _aLez_T_36; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_38 = unsignedAReg[7] ? 5'h18 : _aLez_T_37; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_39 = unsignedAReg[8] ? 5'h17 : _aLez_T_38; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_40 = unsignedAReg[9] ? 5'h16 : _aLez_T_39; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_41 = unsignedAReg[10] ? 5'h15 : _aLez_T_40; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_42 = unsignedAReg[11] ? 5'h14 : _aLez_T_41; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_43 = unsignedAReg[12] ? 5'h13 : _aLez_T_42; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_44 = unsignedAReg[13] ? 5'h12 : _aLez_T_43; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_45 = unsignedAReg[14] ? 5'h11 : _aLez_T_44; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_46 = unsignedAReg[15] ? 5'h10 : _aLez_T_45; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_47 = unsignedAReg[16] ? 5'hf : _aLez_T_46; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_48 = unsignedAReg[17] ? 5'he : _aLez_T_47; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_49 = unsignedAReg[18] ? 5'hd : _aLez_T_48; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_50 = unsignedAReg[19] ? 5'hc : _aLez_T_49; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_51 = unsignedAReg[20] ? 5'hb : _aLez_T_50; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_52 = unsignedAReg[21] ? 5'ha : _aLez_T_51; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_53 = unsignedAReg[22] ? 5'h9 : _aLez_T_52; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_54 = unsignedAReg[23] ? 5'h8 : _aLez_T_53; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_55 = unsignedAReg[24] ? 5'h7 : _aLez_T_54; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_56 = unsignedAReg[25] ? 5'h6 : _aLez_T_55; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_57 = unsignedAReg[26] ? 5'h5 : _aLez_T_56; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_58 = unsignedAReg[27] ? 5'h4 : _aLez_T_57; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_59 = unsignedAReg[28] ? 5'h3 : _aLez_T_58; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_60 = unsignedAReg[29] ? 5'h2 : _aLez_T_59; // @[Mux.scala 47:70]
  wire [4:0] _aLez_T_61 = unsignedAReg[30] ? 5'h1 : _aLez_T_60; // @[Mux.scala 47:70]
  wire [4:0] aLez = unsignedAReg[31] ? 5'h0 : _aLez_T_61; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_32 = unsignedDReg[1] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_33 = unsignedDReg[2] ? 5'h1d : _dLez_T_32; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_34 = unsignedDReg[3] ? 5'h1c : _dLez_T_33; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_35 = unsignedDReg[4] ? 5'h1b : _dLez_T_34; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_36 = unsignedDReg[5] ? 5'h1a : _dLez_T_35; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_37 = unsignedDReg[6] ? 5'h19 : _dLez_T_36; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_38 = unsignedDReg[7] ? 5'h18 : _dLez_T_37; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_39 = unsignedDReg[8] ? 5'h17 : _dLez_T_38; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_40 = unsignedDReg[9] ? 5'h16 : _dLez_T_39; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_41 = unsignedDReg[10] ? 5'h15 : _dLez_T_40; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_42 = unsignedDReg[11] ? 5'h14 : _dLez_T_41; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_43 = unsignedDReg[12] ? 5'h13 : _dLez_T_42; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_44 = unsignedDReg[13] ? 5'h12 : _dLez_T_43; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_45 = unsignedDReg[14] ? 5'h11 : _dLez_T_44; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_46 = unsignedDReg[15] ? 5'h10 : _dLez_T_45; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_47 = unsignedDReg[16] ? 5'hf : _dLez_T_46; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_48 = unsignedDReg[17] ? 5'he : _dLez_T_47; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_49 = unsignedDReg[18] ? 5'hd : _dLez_T_48; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_50 = unsignedDReg[19] ? 5'hc : _dLez_T_49; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_51 = unsignedDReg[20] ? 5'hb : _dLez_T_50; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_52 = unsignedDReg[21] ? 5'ha : _dLez_T_51; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_53 = unsignedDReg[22] ? 5'h9 : _dLez_T_52; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_54 = unsignedDReg[23] ? 5'h8 : _dLez_T_53; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_55 = unsignedDReg[24] ? 5'h7 : _dLez_T_54; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_56 = unsignedDReg[25] ? 5'h6 : _dLez_T_55; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_57 = unsignedDReg[26] ? 5'h5 : _dLez_T_56; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_58 = unsignedDReg[27] ? 5'h4 : _dLez_T_57; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_59 = unsignedDReg[28] ? 5'h3 : _dLez_T_58; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_60 = unsignedDReg[29] ? 5'h2 : _dLez_T_59; // @[Mux.scala 47:70]
  wire [4:0] _dLez_T_61 = unsignedDReg[30] ? 5'h1 : _dLez_T_60; // @[Mux.scala 47:70]
  wire [4:0] dLez = unsignedDReg[31] ? 5'h0 : _dLez_T_61; // @[Mux.scala 47:70]
  wire [4:0] _iter_T_2 = dLez - aLez; // @[IntDivMod.scala 36:41]
  wire [4:0] _iter_T_4 = _iter_T_2 + 5'h1; // @[IntDivMod.scala 36:48]
  wire [4:0] iter = aLez > dLez ? 5'h0 : _iter_T_4; // @[IntDivMod.scala 36:17]
  reg [33:0] aReg; // @[IntDivMod.scala 38:21]
  reg [33:0] dReg; // @[IntDivMod.scala 39:21]
  wire [62:0] _GEN_0 = {{31'd0}, unsignedAReg}; // @[IntDivMod.scala 40:42]
  wire [62:0] _aNorm_T = _GEN_0 << aLez; // @[IntDivMod.scala 40:42]
  wire [33:0] aNorm = {2'h0,_aNorm_T[31:0]}; // @[Cat.scala 31:58]
  wire [62:0] _GEN_1 = {{31'd0}, unsignedDReg}; // @[IntDivMod.scala 41:42]
  wire [62:0] _dNorm_T = _GEN_1 << dLez; // @[IntDivMod.scala 41:42]
  wire [33:0] dNorm = {1'h0,_dNorm_T[31:0],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] _dNegNorm_T = ~unsignedDReg; // @[IntDivMod.scala 42:35]
  wire [31:0] _dNegNorm_T_2 = _dNegNorm_T + 32'h1; // @[IntDivMod.scala 42:59]
  wire [62:0] _GEN_2 = {{31'd0}, _dNegNorm_T_2}; // @[IntDivMod.scala 42:65]
  wire [62:0] _dNegNorm_T_3 = _GEN_2 << dLez; // @[IntDivMod.scala 42:65]
  wire [33:0] dNegNorm = {1'h1,_dNegNorm_T_3[31:0],1'h0}; // @[Cat.scala 31:58]
  wire  _iterReg_T = state == 3'h1; // @[IntDivMod.scala 43:38]
  wire  _zeroQReg_T = unsignedAReg < unsignedDReg; // @[IntDivMod.scala 44:41]
  reg  zeroQReg; // @[Reg.scala 16:16]
  reg [4:0] cnt; // @[IntDivMod.scala 46:20]
  wire [4:0] _cnt_next_T_2 = cnt - 5'h1; // @[IntDivMod.scala 47:42]
  wire [4:0] cnt_next = cnt == 5'h0 ? 5'h0 : _cnt_next_T_2; // @[IntDivMod.scala 47:21]
  reg [31:0] Q; // @[IntDivMod.scala 49:18]
  reg [31:0] QN; // @[IntDivMod.scala 50:19]
  wire  sel_pos = aReg[32:31] == 2'h1; // @[IntDivMod.scala 52:37]
  wire  sel_neg = aReg[32:31] == 2'h2; // @[IntDivMod.scala 53:37]
  wire [34:0] _aShift_T = {aReg, 1'h0}; // @[IntDivMod.scala 55:21]
  wire [33:0] aShift = _aShift_T[33:0]; // @[IntDivMod.scala 55:30]
  wire [33:0] _aNext_T_1 = aShift + dNegNorm; // @[IntDivMod.scala 56:35]
  wire [33:0] _aNext_T_3 = aShift + dNorm; // @[IntDivMod.scala 56:67]
  wire [33:0] _aNext_T_4 = sel_neg ? _aNext_T_3 : aShift; // @[IntDivMod.scala 56:50]
  wire [33:0] aNext = sel_pos ? _aNext_T_1 : _aNext_T_4; // @[IntDivMod.scala 56:18]
  wire  remIsNeg = aReg[33]; // @[IntDivMod.scala 58:27]
  wire [31:0] _commonQReg_T_1 = ~QN; // @[IntDivMod.scala 59:58]
  wire [31:0] _commonQReg_T_3 = Q + _commonQReg_T_1; // @[IntDivMod.scala 59:55]
  wire [31:0] _commonQReg_T_5 = Q - QN; // @[IntDivMod.scala 59:75]
  wire  _commonQReg_T_7 = state == 3'h3; // @[IntDivMod.scala 59:87]
  reg [31:0] commonQReg; // @[Reg.scala 16:16]
  wire [31:0] _recoveryR_T_6 = aReg[32:1] + dReg[32:1]; // @[IntDivMod.scala 60:65]
  wire [31:0] recoveryR = remIsNeg ? _recoveryR_T_6 : aReg[32:1]; // @[IntDivMod.scala 60:22]
  wire [31:0] _commonRReg_T = recoveryR >> dLez; // @[IntDivMod.scala 61:40]
  reg [31:0] commonRReg; // @[Reg.scala 16:16]
  wire [31:0] _signedQ_T = ~commonQReg; // @[IntDivMod.scala 63:32]
  wire [31:0] _signedQ_T_2 = _signedQ_T + 32'h1; // @[IntDivMod.scala 63:54]
  wire [31:0] signedQ = qSignReg ? _signedQ_T_2 : commonQReg; // @[IntDivMod.scala 63:20]
  wire [31:0] _signedR_T = ~commonRReg; // @[IntDivMod.scala 64:32]
  wire [31:0] _signedR_T_2 = _signedR_T + 32'h1; // @[IntDivMod.scala 64:54]
  wire [31:0] signedR = rSignReg ? _signedR_T_2 : commonRReg; // @[IntDivMod.scala 64:20]
  wire [31:0] _specialQ_T_2 = overflowReg ? 32'h80000000 : 32'h0; // @[IntDivMod.scala 65:64]
  wire [31:0] specialQ = divByZeroReg ? 32'hffffffff : _specialQ_T_2; // @[IntDivMod.scala 65:21]
  wire  _specialR_T = divByZeroReg | zeroQReg; // @[IntDivMod.scala 67:34]
  wire [31:0] specialR = divByZeroReg | zeroQReg ? rawAReg : 32'h0; // @[IntDivMod.scala 67:21]
  wire  _io_out_bits_q_T_1 = _specialR_T | overflowReg; // @[IntDivMod.scala 69:46]
  wire  _T = 3'h0 == state; // @[IntDivMod.scala 75:16]
  wire  _T_3 = 3'h1 == state; // @[IntDivMod.scala 75:16]
  wire  _T_5 = 3'h2 == state; // @[IntDivMod.scala 75:16]
  wire [2:0] _GEN_14 = cnt_next != 5'h0 ? 3'h2 : 3'h3; // @[IntDivMod.scala 87:{29,37} 88:26]
  wire  _T_7 = 3'h3 == state; // @[IntDivMod.scala 75:16]
  wire  _T_8 = 3'h4 == state; // @[IntDivMod.scala 75:16]
  wire  _T_9 = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_15 = _T_9 ? 3'h0 : state; // @[IntDivMod.scala 16:22 92:{26,34}]
  wire [2:0] _GEN_16 = 3'h4 == state ? _GEN_15 : state; // @[IntDivMod.scala 75:16 16:22]
  wire [2:0] _GEN_17 = 3'h3 == state ? 3'h4 : _GEN_16; // @[IntDivMod.scala 75:16 90:27]
  wire [31:0] _Q_T_1 = {Q[30:0],sel_pos}; // @[Cat.scala 31:58]
  wire [31:0] _QN_T_1 = {QN[30:0],sel_neg}; // @[Cat.scala 31:58]
  wire [4:0] _GEN_26 = _T_8 ? 5'h0 : cnt; // @[IntDivMod.scala 123:11 96:16 46:20]
  wire [4:0] _GEN_27 = _T_7 ? 5'h0 : _GEN_26; // @[IntDivMod.scala 120:11 96:16]
  assign io_in_ready = state == 3'h0; // @[IntDivMod.scala 72:23]
  assign io_out_valid = state == 3'h4; // @[IntDivMod.scala 71:24]
  assign io_out_bits_q = _specialR_T | overflowReg ? specialQ : signedQ; // @[IntDivMod.scala 69:23]
  assign io_out_bits_r = _io_out_bits_q_T_1 ? specialR : signedR; // @[IntDivMod.scala 70:23]
  always @(posedge clock) begin
    if (reset) begin // @[IntDivMod.scala 16:22]
      state <= 3'h0; // @[IntDivMod.scala 16:22]
    end else if (3'h0 == state) begin // @[IntDivMod.scala 75:16]
      if (_qSignReg_T_1) begin // @[IntDivMod.scala 77:25]
        if (overflow | divByZero) begin // @[IntDivMod.scala 78:36]
          state <= 3'h4; // @[IntDivMod.scala 78:44]
        end else begin
          state <= 3'h1; // @[IntDivMod.scala 79:28]
        end
      end
    end else if (3'h1 == state) begin // @[IntDivMod.scala 75:16]
      if (_zeroQReg_T) begin // @[IntDivMod.scala 83:40]
        state <= 3'h4; // @[IntDivMod.scala 83:48]
      end else begin
        state <= 3'h2; // @[IntDivMod.scala 84:26]
      end
    end else if (3'h2 == state) begin // @[IntDivMod.scala 75:16]
      state <= _GEN_14;
    end else begin
      state <= _GEN_17;
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      qSignReg <= _qSignReg_T; // @[Reg.scala 17:22]
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      rSignReg <= aSign; // @[Reg.scala 17:22]
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      rawAReg <= io_in_bits_a; // @[Reg.scala 17:22]
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      if (aSign) begin // @[IntDivMod.scala 22:22]
        unsignedAReg <= _unsignedA_T_2;
      end else begin
        unsignedAReg <= io_in_bits_a;
      end
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      if (dSign) begin // @[IntDivMod.scala 23:22]
        unsignedDReg <= _unsignedD_T_2;
      end else begin
        unsignedDReg <= io_in_bits_d;
      end
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      overflowReg <= overflow; // @[Reg.scala 17:22]
    end
    if (_qSignReg_T_1) begin // @[Reg.scala 17:18]
      divByZeroReg <= divByZero; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[IntDivMod.scala 38:21]
      aReg <= 34'h0; // @[IntDivMod.scala 38:21]
    end else if (_T) begin // @[IntDivMod.scala 96:16]
      aReg <= 34'h0; // @[IntDivMod.scala 98:12]
    end else if (_T_3) begin // @[IntDivMod.scala 96:16]
      if (!(_zeroQReg_T)) begin // @[IntDivMod.scala 103:40]
        aReg <= aNorm; // @[IntDivMod.scala 106:14]
      end
    end else if (_T_5) begin // @[IntDivMod.scala 96:16]
      aReg <= aNext; // @[IntDivMod.scala 115:12]
    end
    if (reset) begin // @[IntDivMod.scala 39:21]
      dReg <= 34'h0; // @[IntDivMod.scala 39:21]
    end else if (_T) begin // @[IntDivMod.scala 96:16]
      dReg <= 34'h0; // @[IntDivMod.scala 99:12]
    end else if (_T_3) begin // @[IntDivMod.scala 96:16]
      if (!(_zeroQReg_T)) begin // @[IntDivMod.scala 103:40]
        dReg <= dNorm; // @[IntDivMod.scala 107:14]
      end
    end
    if (_iterReg_T) begin // @[Reg.scala 17:18]
      zeroQReg <= _zeroQReg_T; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[IntDivMod.scala 46:20]
      cnt <= 5'h0; // @[IntDivMod.scala 46:20]
    end else if (_T) begin // @[IntDivMod.scala 96:16]
      cnt <= 5'h0; // @[IntDivMod.scala 100:11]
    end else if (_T_3) begin // @[IntDivMod.scala 96:16]
      if (_zeroQReg_T) begin // @[IntDivMod.scala 103:40]
        cnt <= 5'h0; // @[IntDivMod.scala 104:13]
      end else begin
        cnt <= iter; // @[IntDivMod.scala 108:13]
      end
    end else if (_T_5) begin // @[IntDivMod.scala 96:16]
      cnt <= cnt_next; // @[IntDivMod.scala 114:11]
    end else begin
      cnt <= _GEN_27;
    end
    if (reset) begin // @[IntDivMod.scala 49:18]
      Q <= 32'h0; // @[IntDivMod.scala 49:18]
    end else if (!(_T)) begin // @[IntDivMod.scala 96:16]
      if (_T_3) begin // @[IntDivMod.scala 96:16]
        if (!(_zeroQReg_T)) begin // @[IntDivMod.scala 103:40]
          Q <= 32'h0; // @[IntDivMod.scala 109:11]
        end
      end else if (_T_5) begin // @[IntDivMod.scala 96:16]
        Q <= _Q_T_1; // @[IntDivMod.scala 116:9]
      end
    end
    if (reset) begin // @[IntDivMod.scala 50:19]
      QN <= 32'h0; // @[IntDivMod.scala 50:19]
    end else if (!(_T)) begin // @[IntDivMod.scala 96:16]
      if (_T_3) begin // @[IntDivMod.scala 96:16]
        if (!(_zeroQReg_T)) begin // @[IntDivMod.scala 103:40]
          QN <= 32'h0; // @[IntDivMod.scala 110:12]
        end
      end else if (_T_5) begin // @[IntDivMod.scala 96:16]
        QN <= _QN_T_1; // @[IntDivMod.scala 117:10]
      end
    end
    if (_commonQReg_T_7) begin // @[Reg.scala 17:18]
      if (remIsNeg) begin // @[IntDivMod.scala 59:33]
        commonQReg <= _commonQReg_T_3;
      end else begin
        commonQReg <= _commonQReg_T_5;
      end
    end
    if (_commonQReg_T_7) begin // @[Reg.scala 17:18]
      commonRReg <= _commonRReg_T; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  qSignReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  rawAReg = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  unsignedAReg = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  unsignedDReg = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  overflowReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  divByZeroReg = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  aReg = _RAND_8[33:0];
  _RAND_9 = {2{`RANDOM}};
  dReg = _RAND_9[33:0];
  _RAND_10 = {1{`RANDOM}};
  zeroQReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cnt = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  Q = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  QN = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  commonQReg = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  commonRReg = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SrtTable(
  input  [2:0] io_d,
  input  [7:0] io_y,
  output [2:0] io_q
);
  wire  _T_1 = $signed(io_y) >= 8'sh18; // @[util.scala 166:58]
  wire  _T_3 = $signed(io_y) >= 8'sh8; // @[util.scala 166:58]
  wire  _T_5 = $signed(io_y) >= -8'sh8; // @[util.scala 166:58]
  wire  _T_7 = $signed(io_y) >= -8'sh1a; // @[util.scala 166:58]
  wire  _T_9 = $signed(io_y) >= 8'sh1c; // @[util.scala 166:58]
  wire  _T_11 = $signed(io_y) >= -8'sha; // @[util.scala 166:58]
  wire  _T_13 = $signed(io_y) >= -8'sh1c; // @[util.scala 166:58]
  wire  _T_15 = $signed(io_y) >= 8'sh20; // @[util.scala 166:58]
  wire  _T_17 = $signed(io_y) >= -8'shc; // @[util.scala 166:58]
  wire  _T_19 = $signed(io_y) >= -8'sh20; // @[util.scala 166:58]
  wire  _T_21 = $signed(io_y) >= -8'sh22; // @[util.scala 166:58]
  wire  _T_23 = $signed(io_y) >= 8'sh24; // @[util.scala 166:58]
  wire  _T_25 = $signed(io_y) >= 8'shc; // @[util.scala 166:58]
  wire  _T_27 = $signed(io_y) >= -8'sh24; // @[util.scala 166:58]
  wire  _T_29 = $signed(io_y) >= 8'sh28; // @[util.scala 166:58]
  wire  _T_31 = $signed(io_y) >= -8'sh10; // @[util.scala 166:58]
  wire  _T_33 = $signed(io_y) >= -8'sh28; // @[util.scala 166:58]
  wire  _T_35 = $signed(io_y) >= 8'sh10; // @[util.scala 166:58]
  wire  _T_37 = $signed(io_y) >= -8'sh2c; // @[util.scala 166:58]
  wire  _T_39 = $signed(io_y) >= 8'sh30; // @[util.scala 166:58]
  wire  _T_41 = $signed(io_y) >= -8'sh2e; // @[util.scala 166:58]
  wire [2:0] _io_q_T = _T_7 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_1 = _T_5 ? $signed(3'sh0) : $signed(_io_q_T); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_2 = _T_3 ? $signed(3'sh1) : $signed(_io_q_T_1); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_3 = _T_1 ? $signed(3'sh2) : $signed(_io_q_T_2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_4 = _T_13 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_5 = _T_11 ? $signed(3'sh0) : $signed(_io_q_T_4); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_6 = _T_3 ? $signed(3'sh1) : $signed(_io_q_T_5); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_7 = _T_9 ? $signed(3'sh2) : $signed(_io_q_T_6); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_8 = _T_19 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_9 = _T_17 ? $signed(3'sh0) : $signed(_io_q_T_8); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_10 = _T_3 ? $signed(3'sh1) : $signed(_io_q_T_9); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_11 = _T_15 ? $signed(3'sh2) : $signed(_io_q_T_10); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_12 = _T_21 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_13 = _T_17 ? $signed(3'sh0) : $signed(_io_q_T_12); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_14 = _T_3 ? $signed(3'sh1) : $signed(_io_q_T_13); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_15 = _T_15 ? $signed(3'sh2) : $signed(_io_q_T_14); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_16 = _T_27 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_17 = _T_17 ? $signed(3'sh0) : $signed(_io_q_T_16); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_18 = _T_25 ? $signed(3'sh1) : $signed(_io_q_T_17); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_19 = _T_23 ? $signed(3'sh2) : $signed(_io_q_T_18); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_20 = _T_33 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_21 = _T_31 ? $signed(3'sh0) : $signed(_io_q_T_20); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_22 = _T_25 ? $signed(3'sh1) : $signed(_io_q_T_21); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_23 = _T_29 ? $signed(3'sh2) : $signed(_io_q_T_22); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_24 = _T_37 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_25 = _T_31 ? $signed(3'sh0) : $signed(_io_q_T_24); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_26 = _T_35 ? $signed(3'sh1) : $signed(_io_q_T_25); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_27 = _T_29 ? $signed(3'sh2) : $signed(_io_q_T_26); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_28 = _T_41 ? $signed(-3'sh1) : $signed(-3'sh2); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_29 = _T_31 ? $signed(3'sh0) : $signed(_io_q_T_28); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_30 = _T_35 ? $signed(3'sh1) : $signed(_io_q_T_29); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_31 = _T_39 ? $signed(3'sh2) : $signed(_io_q_T_30); // @[Mux.scala 101:16]
  wire [2:0] _io_q_T_33 = 3'h1 == io_d ? $signed(_io_q_T_7) : $signed(_io_q_T_3); // @[Mux.scala 81:58]
  wire [2:0] _io_q_T_35 = 3'h2 == io_d ? $signed(_io_q_T_11) : $signed(_io_q_T_33); // @[Mux.scala 81:58]
  wire [2:0] _io_q_T_37 = 3'h3 == io_d ? $signed(_io_q_T_15) : $signed(_io_q_T_35); // @[Mux.scala 81:58]
  wire [2:0] _io_q_T_39 = 3'h4 == io_d ? $signed(_io_q_T_19) : $signed(_io_q_T_37); // @[Mux.scala 81:58]
  wire [2:0] _io_q_T_41 = 3'h5 == io_d ? $signed(_io_q_T_23) : $signed(_io_q_T_39); // @[Mux.scala 81:58]
  wire [2:0] _io_q_T_43 = 3'h6 == io_d ? $signed(_io_q_T_27) : $signed(_io_q_T_41); // @[Mux.scala 81:58]
  assign io_q = 3'h7 == io_d ? $signed(_io_q_T_31) : $signed(_io_q_T_43); // @[Mux.scala 81:58]
endmodule
module OnTheFlyConv(
  input         clock,
  input         io_resetSqrt,
  input         io_resetDiv,
  input         io_enable,
  input  [2:0]  io_qi,
  output [30:0] io_QM,
  output [30:0] io_Q,
  output [30:0] io_F
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [30:0] Q; // @[util.scala 191:18]
  reg [30:0] QM; // @[util.scala 191:18]
  reg [30:0] mask; // @[util.scala 193:17]
  reg [30:0] b_111; // @[util.scala 194:26]
  reg [30:0] b_1100; // @[util.scala 194:26]
  wire [28:0] _mask_T_2 = mask[30:2]; // @[util.scala 200:18]
  reg [27:0] b_01; // @[util.scala 204:35]
  reg [27:0] b_10; // @[util.scala 204:35]
  reg [27:0] b_11; // @[util.scala 204:35]
  wire [30:0] negQ = ~Q; // @[util.scala 216:14]
  wire [1:0] _T_3 = io_qi[0] ? 2'h1 : 2'h2; // @[util.scala 224:24]
  wire [33:0] _GEN_3 = {{3'd0}, negQ}; // @[util.scala 224:18]
  wire [33:0] _T_4 = _GEN_3 << _T_3; // @[util.scala 224:18]
  wire [30:0] _T_7 = $signed(mask) >>> io_qi[0]; // @[util.scala 224:82]
  wire [33:0] _GEN_18 = {{3'd0}, _T_7}; // @[util.scala 224:55]
  wire [33:0] _T_8 = _T_4 & _GEN_18; // @[util.scala 224:55]
  wire [33:0] _GEN_19 = {{3'd0}, b_111}; // @[util.scala 224:87]
  wire [33:0] _T_9 = _T_8 | _GEN_19; // @[util.scala 224:87]
  wire [33:0] _GEN_21 = {{3'd0}, b_1100}; // @[util.scala 224:87]
  wire [33:0] _T_18 = _T_8 | _GEN_21; // @[util.scala 224:87]
  wire [33:0] _GEN_4 = {{3'd0}, QM}; // @[util.scala 224:18]
  wire [33:0] _T_22 = _GEN_4 << _T_3; // @[util.scala 224:18]
  wire [33:0] _T_26 = _T_22 & _GEN_18; // @[util.scala 224:55]
  wire [33:0] _T_27 = _T_26 | _GEN_19; // @[util.scala 224:87]
  wire [33:0] _T_36 = _T_26 | _GEN_21; // @[util.scala 224:87]
  wire [33:0] _sqrtToCsa_T_2 = 3'h1 == io_qi ? _T_9 : 34'h0; // @[Mux.scala 81:58]
  wire [33:0] _sqrtToCsa_T_4 = 3'h2 == io_qi ? _T_18 : _sqrtToCsa_T_2; // @[Mux.scala 81:58]
  wire [33:0] _sqrtToCsa_T_6 = 3'h7 == io_qi ? _T_27 : _sqrtToCsa_T_4; // @[Mux.scala 81:58]
  wire [33:0] sqrtToCsa = 3'h6 == io_qi ? _T_36 : _sqrtToCsa_T_6; // @[Mux.scala 81:58]
  wire [30:0] _GEN_26 = {{3'd0}, b_01}; // @[util.scala 230:21]
  wire [30:0] Q_load_01 = Q | _GEN_26; // @[util.scala 230:21]
  wire [30:0] _GEN_27 = {{3'd0}, b_10}; // @[util.scala 231:21]
  wire [30:0] Q_load_10 = Q | _GEN_27; // @[util.scala 231:21]
  wire [30:0] QM_load_01 = QM | _GEN_26; // @[util.scala 232:23]
  wire [30:0] QM_load_10 = QM | _GEN_27; // @[util.scala 233:23]
  wire [30:0] _GEN_30 = {{3'd0}, b_11}; // @[util.scala 234:23]
  wire [30:0] QM_load_11 = QM | _GEN_30; // @[util.scala 234:23]
  wire [30:0] _Q_T_3 = 3'h0 == io_qi ? Q : 31'h0; // @[Mux.scala 81:58]
  wire [30:0] _Q_T_5 = 3'h1 == io_qi ? Q_load_01 : _Q_T_3; // @[Mux.scala 81:58]
  wire [30:0] _Q_T_7 = 3'h2 == io_qi ? Q_load_10 : _Q_T_5; // @[Mux.scala 81:58]
  wire [30:0] _Q_T_9 = 3'h7 == io_qi ? QM_load_11 : _Q_T_7; // @[Mux.scala 81:58]
  wire [30:0] _QM_T_2 = 3'h1 == io_qi ? Q : 31'h0; // @[Mux.scala 81:58]
  wire [30:0] _QM_T_4 = 3'h2 == io_qi ? Q_load_01 : _QM_T_2; // @[Mux.scala 81:58]
  wire [30:0] _QM_T_6 = 3'h0 == io_qi ? QM_load_11 : _QM_T_4; // @[Mux.scala 81:58]
  wire [30:0] _QM_T_8 = 3'h7 == io_qi ? QM_load_10 : _QM_T_6; // @[Mux.scala 81:58]
  assign io_QM = QM; // @[util.scala 261:9]
  assign io_Q = Q; // @[util.scala 262:8]
  assign io_F = sqrtToCsa[30:0]; // @[util.scala 260:8]
  always @(posedge clock) begin
    if (io_resetSqrt) begin // @[util.scala 236:21]
      Q <= 31'h10000000; // @[util.scala 237:7]
    end else if (io_resetDiv) begin // @[util.scala 239:26]
      Q <= 31'h0; // @[util.scala 240:7]
    end else if (io_enable) begin // @[util.scala 242:24]
      if (3'h6 == io_qi) begin // @[Mux.scala 81:58]
        Q <= QM_load_10;
      end else begin
        Q <= _Q_T_9;
      end
    end
    if (io_resetSqrt) begin // @[util.scala 236:21]
      QM <= 31'h0; // @[util.scala 238:8]
    end else if (io_resetDiv) begin // @[util.scala 239:26]
      QM <= 31'h0; // @[util.scala 241:8]
    end else if (io_enable) begin // @[util.scala 242:24]
      if (3'h6 == io_qi) begin // @[Mux.scala 81:58]
        QM <= QM_load_01;
      end else begin
        QM <= _QM_T_8;
      end
    end
    if (io_resetSqrt) begin // @[util.scala 195:21]
      mask <= 31'sh40000000; // @[util.scala 196:10]
    end else if (io_enable) begin // @[util.scala 199:24]
      mask <= {{2{_mask_T_2[28]}},_mask_T_2}; // @[util.scala 200:10]
    end
    if (io_resetSqrt) begin // @[util.scala 195:21]
      b_111 <= 31'h1c000000; // @[util.scala 197:11]
    end else if (io_enable) begin // @[util.scala 199:24]
      b_111 <= {{2'd0}, b_111[30:2]}; // @[util.scala 201:11]
    end
    if (io_resetSqrt) begin // @[util.scala 195:21]
      b_1100 <= 31'h30000000; // @[util.scala 198:12]
    end else if (io_enable) begin // @[util.scala 199:24]
      b_1100 <= {{2'd0}, b_1100[30:2]}; // @[util.scala 202:12]
    end
    if (io_resetSqrt | io_resetDiv) begin // @[util.scala 206:36]
      b_01 <= 28'h4000000; // @[util.scala 207:10]
    end else if (io_enable) begin // @[util.scala 210:24]
      b_01 <= {{2'd0}, b_01[27:2]}; // @[util.scala 211:10]
    end
    if (io_resetSqrt | io_resetDiv) begin // @[util.scala 206:36]
      b_10 <= 28'h8000000; // @[util.scala 208:10]
    end else if (io_enable) begin // @[util.scala 210:24]
      b_10 <= {{2'd0}, b_10[27:2]}; // @[util.scala 212:10]
    end
    if (io_resetSqrt | io_resetDiv) begin // @[util.scala 206:36]
      b_11 <= 28'hc000000; // @[util.scala 209:10]
    end else if (io_enable) begin // @[util.scala 210:24]
      b_11 <= {{2'd0}, b_11[27:2]}; // @[util.scala 213:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  Q = _RAND_0[30:0];
  _RAND_1 = {1{`RANDOM}};
  QM = _RAND_1[30:0];
  _RAND_2 = {1{`RANDOM}};
  mask = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  b_111 = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  b_1100 = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  b_01 = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  b_10 = _RAND_6[27:0];
  _RAND_7 = {1{`RANDOM}};
  b_11 = _RAND_7[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSA32(
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  output [31:0] io_out_0,
  output [31:0] io_out_1
);
  wire [31:0] _s_T = io_in_0 ^ io_in_1; // @[util.scala 271:13]
  wire [31:0] _co_T = io_in_0 & io_in_1; // @[util.scala 272:14]
  wire [31:0] _co_T_2 = _s_T & io_in_2; // @[util.scala 272:26]
  assign io_out_0 = _s_T ^ io_in_2; // @[util.scala 271:17]
  assign io_out_1 = _co_T | _co_T_2; // @[util.scala 272:18]
endmodule
module FracDivSqrt(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [27:0] io_in_bits_a,
  input  [27:0] io_in_bits_b,
  input         io_in_bits_isDiv,
  input         io_out_ready,
  output        io_out_valid,
  output [27:0] io_out_bits_quot,
  output        io_out_bits_isZeroRem
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] table__io_d; // @[FloatDivSqrt.scala 45:21]
  wire [7:0] table__io_y; // @[FloatDivSqrt.scala 45:21]
  wire [2:0] table__io_q; // @[FloatDivSqrt.scala 45:21]
  wire  conv_clock; // @[FloatDivSqrt.scala 46:20]
  wire  conv_io_resetSqrt; // @[FloatDivSqrt.scala 46:20]
  wire  conv_io_resetDiv; // @[FloatDivSqrt.scala 46:20]
  wire  conv_io_enable; // @[FloatDivSqrt.scala 46:20]
  wire [2:0] conv_io_qi; // @[FloatDivSqrt.scala 46:20]
  wire [30:0] conv_io_QM; // @[FloatDivSqrt.scala 46:20]
  wire [30:0] conv_io_Q; // @[FloatDivSqrt.scala 46:20]
  wire [30:0] conv_io_F; // @[FloatDivSqrt.scala 46:20]
  wire [31:0] csa_io_in_0; // @[FloatDivSqrt.scala 47:19]
  wire [31:0] csa_io_in_1; // @[FloatDivSqrt.scala 47:19]
  wire [31:0] csa_io_in_2; // @[FloatDivSqrt.scala 47:19]
  wire [31:0] csa_io_out_0; // @[FloatDivSqrt.scala 47:19]
  wire [31:0] csa_io_out_1; // @[FloatDivSqrt.scala 47:19]
  wire  _isDivReg_T = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  reg  isDivReg; // @[Reg.scala 16:16]
  reg [27:0] divisor; // @[Reg.scala 16:16]
  reg [1:0] state; // @[FloatDivSqrt.scala 23:22]
  wire  _cnt_T = state == 2'h0; // @[FloatDivSqrt.scala 25:38]
  wire  _cnt_T_1 = state == 2'h1; // @[FloatDivSqrt.scala 25:56]
  wire  _cnt_T_2 = state == 2'h0 | state == 2'h1; // @[FloatDivSqrt.scala 25:48]
  reg [3:0] cnt; // @[Reg.scala 16:16]
  wire [3:0] _cnt_next_T_2 = cnt - 4'h1; // @[FloatDivSqrt.scala 26:50]
  wire [3:0] cnt_next = _cnt_T ? 4'he : _cnt_next_T_2; // @[FloatDivSqrt.scala 26:18]
  reg  firstCycle; // @[FloatDivSqrt.scala 28:27]
  wire  _T_3 = cnt_next == 4'h0; // @[FloatDivSqrt.scala 35:20]
  wire [1:0] _GEN_5 = io_out_valid ? 2'h0 : state; // @[FloatDivSqrt.scala 23:22 39:{24,32}]
  wire [1:0] _GEN_6 = 2'h3 == state ? _GEN_5 : state; // @[FloatDivSqrt.scala 30:16 23:22]
  reg [31:0] ws; // @[FloatDivSqrt.scala 43:19]
  reg [31:0] wc; // @[FloatDivSqrt.scala 43:19]
  wire [28:0] S = conv_io_Q[30:2]; // @[FloatDivSqrt.scala 50:21]
  wire  s4 = S[22]; // @[FloatDivSqrt.scala 51:66]
  wire  s3 = S[23]; // @[FloatDivSqrt.scala 51:66]
  wire  s2 = S[24]; // @[FloatDivSqrt.scala 51:66]
  wire  s0 = S[26]; // @[FloatDivSqrt.scala 51:66]
  wire [2:0] _sqrt_d_T = {s2,s3,s4}; // @[Cat.scala 31:58]
  wire [2:0] _sqrt_d_T_1 = s0 ? 3'h7 : _sqrt_d_T; // @[FloatDivSqrt.scala 52:50]
  wire [2:0] sqrt_d = firstCycle ? 3'h5 : _sqrt_d_T_1; // @[FloatDivSqrt.scala 52:19]
  wire [2:0] div_d = divisor[26:24]; // @[FloatDivSqrt.scala 53:22]
  wire [7:0] sqrt_y = ws[31:24] + wc[31:24]; // @[FloatDivSqrt.scala 54:33]
  wire [7:0] div_y = ws[30:23] + wc[30:23]; // @[FloatDivSqrt.scala 55:32]
  wire [28:0] _dx2_T = {divisor, 1'h0}; // @[FloatDivSqrt.scala 67:18]
  wire [31:0] dx1 = {{4'd0}, divisor}; // @[FloatDivSqrt.scala 65:40 66:7]
  wire [31:0] neg_dx1 = ~dx1; // @[FloatDivSqrt.scala 68:14]
  wire [32:0] _neg_dx2_T = {neg_dx1, 1'h0}; // @[FloatDivSqrt.scala 69:22]
  wire [31:0] _divCsaIn_T_6 = 3'h7 == table__io_q ? dx1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] dx2 = {{3'd0}, _dx2_T}; // @[FloatDivSqrt.scala 65:40 67:7]
  wire [31:0] _divCsaIn_T_8 = 3'h6 == table__io_q ? dx2 : _divCsaIn_T_6; // @[Mux.scala 81:58]
  wire [31:0] _divCsaIn_T_10 = 3'h1 == table__io_q ? neg_dx1 : _divCsaIn_T_8; // @[Mux.scala 81:58]
  wire [31:0] neg_dx2 = _neg_dx2_T[31:0]; // @[FloatDivSqrt.scala 65:40 69:11]
  wire [31:0] divCsaIn = 3'h2 == table__io_q ? neg_dx2 : _divCsaIn_T_10; // @[Mux.scala 81:58]
  wire [31:0] _GEN_16 = {{30'd0}, table__io_q[1:0]}; // @[FloatDivSqrt.scala 79:52]
  wire [31:0] _csa_io_in_1_T_4 = wc | _GEN_16; // @[FloatDivSqrt.scala 79:52]
  wire [29:0] _sqrtWsInit_T = {2'h0,io_in_bits_a}; // @[Cat.scala 31:58]
  wire [29:0] _sqrtWsInit_T_3 = _sqrtWsInit_T - 30'h10000000; // @[FloatDivSqrt.scala 84:42]
  wire [31:0] sqrtWsInit = {_sqrtWsInit_T_3,2'h0}; // @[Cat.scala 31:58]
  wire [31:0] _ws_T = io_in_bits_isDiv ? {{4'd0}, io_in_bits_a} : sqrtWsInit; // @[FloatDivSqrt.scala 88:14]
  wire [33:0] _ws_T_2 = {csa_io_out_0, 2'h0}; // @[FloatDivSqrt.scala 91:59]
  wire [33:0] _ws_T_3 = _T_3 ? {{2'd0}, csa_io_out_0} : _ws_T_2; // @[FloatDivSqrt.scala 91:14]
  wire [32:0] _wc_T_1 = {csa_io_out_1, 1'h0}; // @[FloatDivSqrt.scala 92:44]
  wire [34:0] _wc_T_2 = {csa_io_out_1, 3'h0}; // @[FloatDivSqrt.scala 92:62]
  wire [34:0] _wc_T_3 = _T_3 ? {{2'd0}, _wc_T_1} : _wc_T_2; // @[FloatDivSqrt.scala 92:14]
  wire [33:0] _GEN_10 = _cnt_T_1 ? _ws_T_3 : {{2'd0}, ws}; // @[FloatDivSqrt.scala 43:19 90:35 91:8]
  wire [34:0] _GEN_11 = _cnt_T_1 ? _wc_T_3 : {{3'd0}, wc}; // @[FloatDivSqrt.scala 43:19 90:35 92:8]
  wire [33:0] _GEN_12 = _isDivReg_T ? {{2'd0}, _ws_T} : _GEN_10; // @[FloatDivSqrt.scala 87:21 88:8]
  wire [34:0] _GEN_13 = _isDivReg_T ? 35'h0 : _GEN_11; // @[FloatDivSqrt.scala 87:21 89:8]
  wire [31:0] rem = ws + wc; // @[FloatDivSqrt.scala 94:16]
  wire  _remSignReg_T_2 = state == 2'h2; // @[FloatDivSqrt.scala 95:57]
  reg  remSignReg; // @[Reg.scala 16:16]
  wire  _isZeroRemReg_T = rem == 32'h0; // @[FloatDivSqrt.scala 96:35]
  reg  isZeroRemReg; // @[Reg.scala 16:16]
  wire [30:0] _io_out_bits_quot_T = remSignReg ? conv_io_QM : conv_io_Q; // @[FloatDivSqrt.scala 99:26]
  wire [30:0] _io_out_bits_quot_T_2 = _io_out_bits_quot_T >> ~isDivReg; // @[FloatDivSqrt.scala 99:62]
  SrtTable table_ ( // @[FloatDivSqrt.scala 45:21]
    .io_d(table__io_d),
    .io_y(table__io_y),
    .io_q(table__io_q)
  );
  OnTheFlyConv conv ( // @[FloatDivSqrt.scala 46:20]
    .clock(conv_clock),
    .io_resetSqrt(conv_io_resetSqrt),
    .io_resetDiv(conv_io_resetDiv),
    .io_enable(conv_io_enable),
    .io_qi(conv_io_qi),
    .io_QM(conv_io_QM),
    .io_Q(conv_io_Q),
    .io_F(conv_io_F)
  );
  CSA32 csa ( // @[FloatDivSqrt.scala 47:19]
    .io_in_0(csa_io_in_0),
    .io_in_1(csa_io_in_1),
    .io_in_2(csa_io_in_2),
    .io_out_0(csa_io_out_0),
    .io_out_1(csa_io_out_1)
  );
  assign io_in_ready = state == 2'h0; // @[FloatDivSqrt.scala 97:24]
  assign io_out_valid = state == 2'h3; // @[FloatDivSqrt.scala 98:25]
  assign io_out_bits_quot = _io_out_bits_quot_T_2[27:0]; // @[FloatDivSqrt.scala 99:20]
  assign io_out_bits_isZeroRem = isZeroRemReg; // @[FloatDivSqrt.scala 100:25]
  assign table__io_d = isDivReg ? div_d : sqrt_d; // @[FloatDivSqrt.scala 57:20]
  assign table__io_y = isDivReg ? div_y : sqrt_y; // @[FloatDivSqrt.scala 58:20]
  assign conv_clock = clock;
  assign conv_io_resetSqrt = _isDivReg_T & ~io_in_bits_isDiv; // @[FloatDivSqrt.scala 60:35]
  assign conv_io_resetDiv = _isDivReg_T & io_in_bits_isDiv; // @[FloatDivSqrt.scala 61:34]
  assign conv_io_enable = state == 2'h1; // @[FloatDivSqrt.scala 62:26]
  assign conv_io_qi = table__io_q; // @[FloatDivSqrt.scala 63:14]
  assign csa_io_in_0 = ws; // @[FloatDivSqrt.scala 78:16]
  assign csa_io_in_1 = isDivReg & ~table__io_q[2] ? _csa_io_in_1_T_4 : wc; // @[FloatDivSqrt.scala 79:22]
  assign csa_io_in_2 = isDivReg ? divCsaIn : {{1'd0}, conv_io_F}; // @[FloatDivSqrt.scala 80:22]
  always @(posedge clock) begin
    if (_isDivReg_T) begin // @[Reg.scala 17:18]
      isDivReg <= io_in_bits_isDiv; // @[Reg.scala 17:22]
    end
    if (_isDivReg_T) begin // @[Reg.scala 17:18]
      divisor <= io_in_bits_b; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FloatDivSqrt.scala 23:22]
      state <= 2'h0; // @[FloatDivSqrt.scala 23:22]
    end else if (2'h0 == state) begin // @[FloatDivSqrt.scala 30:16]
      if (_isDivReg_T) begin // @[FloatDivSqrt.scala 32:23]
        state <= 2'h1; // @[FloatDivSqrt.scala 32:31]
      end
    end else if (2'h1 == state) begin // @[FloatDivSqrt.scala 30:16]
      if (cnt_next == 4'h0) begin // @[FloatDivSqrt.scala 35:27]
        state <= 2'h2; // @[FloatDivSqrt.scala 35:35]
      end
    end else if (2'h2 == state) begin // @[FloatDivSqrt.scala 30:16]
      state <= 2'h3; // @[FloatDivSqrt.scala 37:27]
    end else begin
      state <= _GEN_6;
    end
    if (_cnt_T_2) begin // @[Reg.scala 17:18]
      if (_cnt_T) begin // @[FloatDivSqrt.scala 26:18]
        cnt <= 4'he;
      end else begin
        cnt <= _cnt_next_T_2;
      end
    end
    firstCycle <= io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
    ws <= _GEN_12[31:0];
    wc <= _GEN_13[31:0];
    if (_remSignReg_T_2) begin // @[Reg.scala 17:18]
      remSignReg <= rem[31]; // @[Reg.scala 17:22]
    end
    if (_remSignReg_T_2) begin // @[Reg.scala 17:18]
      isZeroRemReg <= _isZeroRemReg_T; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isDivReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  divisor = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  cnt = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  firstCycle = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ws = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  wc = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  remSignReg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  isZeroRemReg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FloatDivSqrt(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_op,
  input  [31:0] io_in_bits_a,
  input  [31:0] io_in_bits_b,
  input  [2:0]  io_in_bits_rm,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] classify_a_io_in; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isNegInf; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isNegNormal; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isNegSubnormal; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isNegZero; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isPosZero; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isPosSubnormal; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isPosNormal; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isPosInf; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isSNaN; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isQNaN; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isNaN; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isInf; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isInfOrNaN; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isSubnormal; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isZero; // @[FloatDivSqrt.scala 119:26]
  wire  classify_a_io_isSubnormalOrZero; // @[FloatDivSqrt.scala 119:26]
  wire [31:0] classify_b_io_in; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isNegInf; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isNegNormal; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isNegSubnormal; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isNegZero; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isPosZero; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isPosSubnormal; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isPosNormal; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isPosInf; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isSNaN; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isQNaN; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isNaN; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isInf; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isInfOrNaN; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isSubnormal; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isZero; // @[FloatDivSqrt.scala 122:26]
  wire  classify_b_io_isSubnormalOrZero; // @[FloatDivSqrt.scala 122:26]
  wire  fracDivSqrt_clock; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_reset; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_io_in_ready; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_io_in_valid; // @[FloatDivSqrt.scala 205:27]
  wire [27:0] fracDivSqrt_io_in_bits_a; // @[FloatDivSqrt.scala 205:27]
  wire [27:0] fracDivSqrt_io_in_bits_b; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_io_in_bits_isDiv; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_io_out_ready; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_io_out_valid; // @[FloatDivSqrt.scala 205:27]
  wire [27:0] fracDivSqrt_io_out_bits_quot; // @[FloatDivSqrt.scala 205:27]
  wire  fracDivSqrt_io_out_bits_isZeroRem; // @[FloatDivSqrt.scala 205:27]
  wire [2:0] rounding_io_in_rm; // @[FloatDivSqrt.scala 237:24]
  wire [23:0] rounding_io_in_frac; // @[FloatDivSqrt.scala 237:24]
  wire  rounding_io_in_sign; // @[FloatDivSqrt.scala 237:24]
  wire  rounding_io_in_guard; // @[FloatDivSqrt.scala 237:24]
  wire  rounding_io_in_round; // @[FloatDivSqrt.scala 237:24]
  wire  rounding_io_in_sticky; // @[FloatDivSqrt.scala 237:24]
  wire [23:0] rounding_io_out_fracRounded; // @[FloatDivSqrt.scala 237:24]
  wire  rounding_io_out_fracCout; // @[FloatDivSqrt.scala 237:24]
  reg [2:0] state; // @[FloatDivSqrt.scala 110:22]
  wire  _rmReg_T = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  reg [2:0] rmReg; // @[Reg.scala 16:16]
  wire  isDiv = io_in_bits_op == 3'h0; // @[FloatDivSqrt.scala 114:28]
  reg  isDivReg; // @[Reg.scala 16:16]
  wire [22:0] f32_frac = io_in_bits_a[22:0]; // @[util.scala 46:46]
  wire [7:0] f32_exp = io_in_bits_a[30:23]; // @[util.scala 46:46]
  wire  f32_sign = io_in_bits_a[31]; // @[util.scala 46:46]
  wire [8:0] _exp_T = {1'h0,f32_exp}; // @[Cat.scala 31:58]
  wire  _fracExt_T = ~classify_a_io_isSubnormalOrZero; // @[FloatDivSqrt.scala 129:23]
  wire [23:0] aFrac = {_fracExt_T,f32_frac}; // @[Cat.scala 31:58]
  wire [8:0] aExp = _exp_T - 9'h7f; // @[FloatDivSqrt.scala 130:20]
  wire [22:0] f32_1_frac = io_in_bits_b[22:0]; // @[util.scala 46:46]
  wire [7:0] f32_1_exp = io_in_bits_b[30:23]; // @[util.scala 46:46]
  wire  f32_1_sign = io_in_bits_b[31]; // @[util.scala 46:46]
  wire [8:0] _exp_T_3 = {1'h0,f32_1_exp}; // @[Cat.scala 31:58]
  wire  _fracExt_T_1 = ~classify_b_io_isSubnormalOrZero; // @[FloatDivSqrt.scala 129:23]
  wire [23:0] bFrac = {_fracExt_T_1,f32_1_frac}; // @[Cat.scala 31:58]
  wire [8:0] bExp = _exp_T_3 - 9'h7f; // @[FloatDivSqrt.scala 130:20]
  wire  resSign = f32_sign ^ f32_1_sign; // @[FloatDivSqrt.scala 135:23]
  reg  resSignReg; // @[Reg.scala 16:16]
  reg [9:0] aExpReg; // @[FloatDivSqrt.scala 137:20]
  reg [23:0] aFracReg; // @[FloatDivSqrt.scala 138:21]
  wire  aIsOddExp = aExpReg[0]; // @[FloatDivSqrt.scala 139:26]
  reg [9:0] bExpReg; // @[FloatDivSqrt.scala 140:20]
  reg [23:0] bFracReg; // @[FloatDivSqrt.scala 141:21]
  reg  aIsSubnormalReg; // @[Reg.scala 16:16]
  reg  bIsSubnormalReg; // @[Reg.scala 16:16]
  wire  hasNaN = classify_a_io_isNaN | classify_b_io_isNaN; // @[FloatDivSqrt.scala 163:23]
  wire  bothZero = classify_a_io_isZero & classify_b_io_isZero; // @[FloatDivSqrt.scala 164:26]
  wire  bothInf = classify_a_io_isInf & classify_b_io_isInf; // @[FloatDivSqrt.scala 165:24]
  wire  _sqrtInvalid_T_5 = ~isDiv; // @[FloatDivSqrt.scala 167:68]
  wire  sqrtSpecial = (f32_sign | classify_a_io_isInfOrNaN | classify_a_io_isZero) & _sqrtInvalid_T_5; // @[FloatDivSqrt.scala 168:55]
  wire  divInvalid = (bothZero | classify_a_io_isSNaN | classify_b_io_isSNaN | bothInf) & isDiv; // @[FloatDivSqrt.scala 170:64]
  wire  divSpecial = (classify_a_io_isZero | classify_b_io_isZero | hasNaN | classify_b_io_isInf | classify_a_io_isInf)
     & isDiv; // @[FloatDivSqrt.scala 172:71]
  wire  _divSpecialResSel_T = divInvalid | hasNaN; // @[FloatDivSqrt.scala 178:17]
  wire  _divSpecialResSel_T_1 = classify_a_io_isZero | classify_b_io_isInf; // @[FloatDivSqrt.scala 180:14]
  wire [2:0] _divSpecialResSel_T_2 = _divSpecialResSel_T_1 ? 3'h2 : 3'h1; // @[Mux.scala 47:70]
  wire [2:0] _divSpecialResSel_T_3 = classify_b_io_isZero ? 3'h1 : _divSpecialResSel_T_2; // @[Mux.scala 47:70]
  wire [2:0] divSpecialResSel = _divSpecialResSel_T ? 3'h4 : _divSpecialResSel_T_3; // @[Mux.scala 47:70]
  wire [2:0] _sqrtSpecialResSel_T = classify_a_io_isPosInf ? 3'h1 : 3'h4; // @[Mux.scala 101:16]
  wire [2:0] sqrtSpecialResSel = classify_a_io_isZero ? 3'h2 : _sqrtSpecialResSel_T; // @[Mux.scala 101:16]
  wire  specialCase = divSpecial | sqrtSpecial; // @[FloatDivSqrt.scala 187:32]
  reg  specialCaseReg; // @[Reg.scala 16:16]
  wire [2:0] specialResSel = sqrtSpecial ? sqrtSpecialResSel : divSpecialResSel; // @[FloatDivSqrt.scala 189:26]
  wire  sel_Zero = specialResSel[1]; // @[FloatDivSqrt.scala 190:68]
  wire  sel_NaN = specialResSel[2]; // @[FloatDivSqrt.scala 190:68]
  wire [31:0] _specialResult_T_3 = {resSign,31'h0}; // @[Cat.scala 31:58]
  wire [31:0] _specialResult_T_7 = {resSign,31'h7f800000}; // @[Cat.scala 31:58]
  reg [31:0] specialResult; // @[Reg.scala 16:16]
  wire [4:0] _aFracLEZ_T_24 = aFracReg[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_25 = aFracReg[2] ? 5'h14 : _aFracLEZ_T_24; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_26 = aFracReg[3] ? 5'h13 : _aFracLEZ_T_25; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_27 = aFracReg[4] ? 5'h12 : _aFracLEZ_T_26; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_28 = aFracReg[5] ? 5'h11 : _aFracLEZ_T_27; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_29 = aFracReg[6] ? 5'h10 : _aFracLEZ_T_28; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_30 = aFracReg[7] ? 5'hf : _aFracLEZ_T_29; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_31 = aFracReg[8] ? 5'he : _aFracLEZ_T_30; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_32 = aFracReg[9] ? 5'hd : _aFracLEZ_T_31; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_33 = aFracReg[10] ? 5'hc : _aFracLEZ_T_32; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_34 = aFracReg[11] ? 5'hb : _aFracLEZ_T_33; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_35 = aFracReg[12] ? 5'ha : _aFracLEZ_T_34; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_36 = aFracReg[13] ? 5'h9 : _aFracLEZ_T_35; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_37 = aFracReg[14] ? 5'h8 : _aFracLEZ_T_36; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_38 = aFracReg[15] ? 5'h7 : _aFracLEZ_T_37; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_39 = aFracReg[16] ? 5'h6 : _aFracLEZ_T_38; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_40 = aFracReg[17] ? 5'h5 : _aFracLEZ_T_39; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_41 = aFracReg[18] ? 5'h4 : _aFracLEZ_T_40; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_42 = aFracReg[19] ? 5'h3 : _aFracLEZ_T_41; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_43 = aFracReg[20] ? 5'h2 : _aFracLEZ_T_42; // @[Mux.scala 47:70]
  wire [4:0] _aFracLEZ_T_44 = aFracReg[21] ? 5'h1 : _aFracLEZ_T_43; // @[Mux.scala 47:70]
  wire [4:0] aFracLEZ = aFracReg[22] ? 5'h0 : _aFracLEZ_T_44; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_24 = bFracReg[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_25 = bFracReg[2] ? 5'h14 : _bFracLEZ_T_24; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_26 = bFracReg[3] ? 5'h13 : _bFracLEZ_T_25; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_27 = bFracReg[4] ? 5'h12 : _bFracLEZ_T_26; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_28 = bFracReg[5] ? 5'h11 : _bFracLEZ_T_27; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_29 = bFracReg[6] ? 5'h10 : _bFracLEZ_T_28; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_30 = bFracReg[7] ? 5'hf : _bFracLEZ_T_29; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_31 = bFracReg[8] ? 5'he : _bFracLEZ_T_30; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_32 = bFracReg[9] ? 5'hd : _bFracLEZ_T_31; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_33 = bFracReg[10] ? 5'hc : _bFracLEZ_T_32; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_34 = bFracReg[11] ? 5'hb : _bFracLEZ_T_33; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_35 = bFracReg[12] ? 5'ha : _bFracLEZ_T_34; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_36 = bFracReg[13] ? 5'h9 : _bFracLEZ_T_35; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_37 = bFracReg[14] ? 5'h8 : _bFracLEZ_T_36; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_38 = bFracReg[15] ? 5'h7 : _bFracLEZ_T_37; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_39 = bFracReg[16] ? 5'h6 : _bFracLEZ_T_38; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_40 = bFracReg[17] ? 5'h5 : _bFracLEZ_T_39; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_41 = bFracReg[18] ? 5'h4 : _bFracLEZ_T_40; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_42 = bFracReg[19] ? 5'h3 : _bFracLEZ_T_41; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_43 = bFracReg[20] ? 5'h2 : _bFracLEZ_T_42; // @[Mux.scala 47:70]
  wire [4:0] _bFracLEZ_T_44 = bFracReg[21] ? 5'h1 : _bFracLEZ_T_43; // @[Mux.scala 47:70]
  wire [4:0] bFracLEZ = bFracReg[22] ? 5'h0 : _bFracLEZ_T_44; // @[Mux.scala 47:70]
  wire [27:0] _fracDivSqrt_io_in_bits_a_T_1 = {aFracReg,4'h0}; // @[Cat.scala 31:58]
  wire [27:0] _fracDivSqrt_io_in_bits_a_T_2 = {1'h0,aFracReg,3'h0}; // @[Cat.scala 31:58]
  wire  needNormalize = ~fracDivSqrt_io_out_bits_quot[26]; // @[FloatDivSqrt.scala 220:23]
  wire [28:0] _fracNorm_T = {fracDivSqrt_io_out_bits_quot, 1'h0}; // @[FloatDivSqrt.scala 221:54]
  wire [28:0] _fracNorm_T_1 = needNormalize ? _fracNorm_T : {{1'd0}, fracDivSqrt_io_out_bits_quot}; // @[FloatDivSqrt.scala 221:21]
  wire [26:0] fracNorm = _fracNorm_T_1[26:0]; // @[FloatDivSqrt.scala 221:77]
  wire [1:0] _expNorm_T_2 = needNormalize ? 2'h2 : 2'h1; // @[FloatDivSqrt.scala 222:85]
  wire [1:0] _expNorm_T_3 = isDivReg ? {{1'd0}, needNormalize} : _expNorm_T_2; // @[FloatDivSqrt.scala 222:41]
  wire [9:0] _GEN_51 = {{8'd0}, _expNorm_T_3}; // @[FloatDivSqrt.scala 222:36]
  wire [9:0] expNorm = aExpReg - _GEN_51; // @[FloatDivSqrt.scala 222:120]
  wire [9:0] denormShift = -10'sh7e - $signed(expNorm); // @[FloatDivSqrt.scala 224:47]
  wire  _denormShiftReg_T = fracDivSqrt_io_out_ready & fracDivSqrt_io_out_valid; // @[Decoupled.scala 50:35]
  wire [9:0] _fracShifted_T_2 = -10'sh7e - $signed(expNorm); // @[FloatDivSqrt.scala 226:102]
  wire [9:0] _fracShifted_T_3 = denormShift[9] ? 10'h0 : _fracShifted_T_2; // @[FloatDivSqrt.scala 226:48]
  wire [4:0] fracShifted_realShiftAmt = _fracShifted_T_3 > 10'h1a ? 5'h1b : _fracShifted_T_3[4:0]; // @[util.scala 125:27]
  wire [4:0] _fracShifted_mask_T_2 = 5'h1b - fracShifted_realShiftAmt; // @[util.scala 129:48]
  wire [26:0] fracShifted_mask = 27'h7ffffff >> _fracShifted_mask_T_2; // @[util.scala 129:41]
  wire [26:0] fracShifted_x_shifted = fracNorm >> fracShifted_realShiftAmt; // @[util.scala 131:24]
  wire [26:0] _fracShifted_T_5 = fracShifted_mask & fracNorm; // @[util.scala 132:32]
  wire [26:0] _GEN_52 = {{26'd0}, |_fracShifted_T_5}; // @[util.scala 132:23]
  wire [26:0] fracShifted = fracShifted_x_shifted | _GEN_52; // @[util.scala 132:23]
  wire [23:0] fracPostNorm = fracShifted[26:3]; // @[FloatDivSqrt.scala 228:38]
  reg  gReg; // @[FloatDivSqrt.scala 232:21]
  reg  rReg; // @[FloatDivSqrt.scala 233:21]
  reg  sReg; // @[FloatDivSqrt.scala 234:21]
  wire  fracCout = ~aFracReg[23] ? rounding_io_out_fracRounded[23] : rounding_io_out_fracCout; // @[FloatDivSqrt.scala 247:21]
  wire [24:0] _isZeroResult_T = {fracCout,rounding_io_out_fracRounded}; // @[Cat.scala 31:58]
  wire  isZeroResult = ~(|_isZeroResult_T); // @[FloatDivSqrt.scala 251:22]
  wire [9:0] _expRounded_T_7 = $signed(aExpReg) + 10'sh7f; // @[FloatDivSqrt.scala 254:13]
  wire [9:0] _expRounded_T_8 = $signed(denormShift) > 10'sh0 | isZeroResult ? $signed(10'sh0) : $signed(_expRounded_T_7)
    ; // @[FloatDivSqrt.scala 252:23]
  wire [1:0] _expRounded_T_10 = {1'h0,fracCout}; // @[util.scala 76:47]
  wire [9:0] _GEN_53 = {{8{_expRounded_T_10[1]}},_expRounded_T_10}; // @[FloatDivSqrt.scala 255:5]
  wire [9:0] expRounded = $signed(_expRounded_T_8) + $signed(_GEN_53); // @[FloatDivSqrt.scala 255:5]
  wire  _T = 3'h0 == state; // @[FloatDivSqrt.scala 275:16]
  wire [2:0] _GEN_16 = classify_a_io_isSubnormal | classify_b_io_isSubnormal ? 3'h1 : 3'h2; // @[FloatDivSqrt.scala 280:49 281:17 283:16]
  wire  _T_4 = 3'h1 == state; // @[FloatDivSqrt.scala 275:16]
  wire  _T_5 = 3'h2 == state; // @[FloatDivSqrt.scala 275:16]
  wire  _T_6 = 3'h3 == state; // @[FloatDivSqrt.scala 275:16]
  wire [2:0] _GEN_19 = _denormShiftReg_T ? 3'h4 : state; // @[FloatDivSqrt.scala 110:22 290:{38,46}]
  wire  _T_8 = 3'h4 == state; // @[FloatDivSqrt.scala 275:16]
  wire  _T_10 = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_20 = _T_10 ? 3'h0 : state; // @[FloatDivSqrt.scala 110:22 293:{39,46}]
  wire [2:0] _GEN_21 = 3'h5 == state ? _GEN_20 : state; // @[FloatDivSqrt.scala 275:16 110:22]
  wire [2:0] _GEN_22 = 3'h4 == state ? 3'h5 : _GEN_21; // @[FloatDivSqrt.scala 275:16 292:24]
  wire [2:0] _GEN_23 = 3'h3 == state ? _GEN_19 : _GEN_22; // @[FloatDivSqrt.scala 275:16]
  wire [23:0] _GEN_28 = _rmReg_T ? aFrac : aFracReg; // @[FloatDivSqrt.scala 298:25 300:18 138:21]
  wire [23:0] _GEN_30 = _rmReg_T ? bFrac : bFracReg; // @[FloatDivSqrt.scala 298:25 302:18 141:21]
  wire [9:0] _GEN_55 = {{5'd0}, aFracLEZ}; // @[FloatDivSqrt.scala 307:38]
  wire [9:0] _aExpReg_T_3 = aExpReg - _GEN_55; // @[FloatDivSqrt.scala 307:56]
  wire [54:0] _GEN_0 = {{31'd0}, aFracReg}; // @[FloatDivSqrt.scala 308:31]
  wire [54:0] _aFracReg_T = _GEN_0 << aFracLEZ; // @[FloatDivSqrt.scala 308:31]
  wire [55:0] _aFracReg_T_1 = {_aFracReg_T, 1'h0}; // @[FloatDivSqrt.scala 308:44]
  wire [55:0] _GEN_32 = aIsSubnormalReg ? _aFracReg_T_1 : {{32'd0}, aFracReg}; // @[FloatDivSqrt.scala 306:28 308:18 138:21]
  wire [9:0] _GEN_56 = {{5'd0}, bFracLEZ}; // @[FloatDivSqrt.scala 311:38]
  wire [9:0] _bExpReg_T_3 = bExpReg - _GEN_56; // @[FloatDivSqrt.scala 311:56]
  wire [54:0] _GEN_1 = {{31'd0}, bFracReg}; // @[FloatDivSqrt.scala 312:31]
  wire [54:0] _bFracReg_T = _GEN_1 << bFracLEZ; // @[FloatDivSqrt.scala 312:31]
  wire [55:0] _bFracReg_T_1 = {_bFracReg_T, 1'h0}; // @[FloatDivSqrt.scala 312:44]
  wire [55:0] _GEN_34 = bIsSubnormalReg ? _bFracReg_T_1 : {{32'd0}, bFracReg}; // @[FloatDivSqrt.scala 310:28 312:18 141:21]
  wire [9:0] _aExpReg_T_6 = $signed(aExpReg) - $signed(bExpReg); // @[FloatDivSqrt.scala 316:40]
  wire [8:0] _aExpReg_T_7 = aExpReg[9:1]; // @[FloatDivSqrt.scala 316:59]
  wire [8:0] _aExpReg_T_10 = $signed(_aExpReg_T_7) + 9'sh1; // @[FloatDivSqrt.scala 316:72]
  wire [9:0] _GEN_35 = _denormShiftReg_T ? $signed(expNorm) : $signed(aExpReg); // @[FloatDivSqrt.scala 319:38 320:17 137:20]
  wire [23:0] _GEN_36 = _denormShiftReg_T ? fracPostNorm : aFracReg; // @[FloatDivSqrt.scala 319:38 321:18 138:21]
  wire [9:0] _GEN_37 = _T_8 ? $signed(expRounded) : $signed(aExpReg); // @[FloatDivSqrt.scala 296:16 325:15 137:20]
  wire [23:0] _GEN_38 = _T_8 ? rounding_io_out_fracRounded : aFracReg; // @[FloatDivSqrt.scala 296:16 326:16 138:21]
  wire [23:0] _GEN_40 = _T_6 ? _GEN_36 : _GEN_38; // @[FloatDivSqrt.scala 296:16]
  wire [23:0] _GEN_42 = _T_5 ? aFracReg : _GEN_40; // @[FloatDivSqrt.scala 296:16 138:21]
  wire [55:0] _GEN_44 = _T_4 ? _GEN_32 : {{32'd0}, _GEN_42}; // @[FloatDivSqrt.scala 296:16]
  wire [55:0] _GEN_46 = _T_4 ? _GEN_34 : {{32'd0}, bFracReg}; // @[FloatDivSqrt.scala 296:16 141:21]
  wire [55:0] _GEN_48 = _T ? {{32'd0}, _GEN_28} : _GEN_44; // @[FloatDivSqrt.scala 296:16]
  wire [55:0] _GEN_50 = _T ? {{32'd0}, _GEN_30} : _GEN_46; // @[FloatDivSqrt.scala 296:16]
  wire [31:0] commonResult = {resSignReg,aExpReg[7:0],aFracReg[22:0]}; // @[Cat.scala 31:58]
  Classify classify_a ( // @[FloatDivSqrt.scala 119:26]
    .io_in(classify_a_io_in),
    .io_isNegInf(classify_a_io_isNegInf),
    .io_isNegNormal(classify_a_io_isNegNormal),
    .io_isNegSubnormal(classify_a_io_isNegSubnormal),
    .io_isNegZero(classify_a_io_isNegZero),
    .io_isPosZero(classify_a_io_isPosZero),
    .io_isPosSubnormal(classify_a_io_isPosSubnormal),
    .io_isPosNormal(classify_a_io_isPosNormal),
    .io_isPosInf(classify_a_io_isPosInf),
    .io_isSNaN(classify_a_io_isSNaN),
    .io_isQNaN(classify_a_io_isQNaN),
    .io_isNaN(classify_a_io_isNaN),
    .io_isInf(classify_a_io_isInf),
    .io_isInfOrNaN(classify_a_io_isInfOrNaN),
    .io_isSubnormal(classify_a_io_isSubnormal),
    .io_isZero(classify_a_io_isZero),
    .io_isSubnormalOrZero(classify_a_io_isSubnormalOrZero)
  );
  Classify classify_b ( // @[FloatDivSqrt.scala 122:26]
    .io_in(classify_b_io_in),
    .io_isNegInf(classify_b_io_isNegInf),
    .io_isNegNormal(classify_b_io_isNegNormal),
    .io_isNegSubnormal(classify_b_io_isNegSubnormal),
    .io_isNegZero(classify_b_io_isNegZero),
    .io_isPosZero(classify_b_io_isPosZero),
    .io_isPosSubnormal(classify_b_io_isPosSubnormal),
    .io_isPosNormal(classify_b_io_isPosNormal),
    .io_isPosInf(classify_b_io_isPosInf),
    .io_isSNaN(classify_b_io_isSNaN),
    .io_isQNaN(classify_b_io_isQNaN),
    .io_isNaN(classify_b_io_isNaN),
    .io_isInf(classify_b_io_isInf),
    .io_isInfOrNaN(classify_b_io_isInfOrNaN),
    .io_isSubnormal(classify_b_io_isSubnormal),
    .io_isZero(classify_b_io_isZero),
    .io_isSubnormalOrZero(classify_b_io_isSubnormalOrZero)
  );
  FracDivSqrt fracDivSqrt ( // @[FloatDivSqrt.scala 205:27]
    .clock(fracDivSqrt_clock),
    .reset(fracDivSqrt_reset),
    .io_in_ready(fracDivSqrt_io_in_ready),
    .io_in_valid(fracDivSqrt_io_in_valid),
    .io_in_bits_a(fracDivSqrt_io_in_bits_a),
    .io_in_bits_b(fracDivSqrt_io_in_bits_b),
    .io_in_bits_isDiv(fracDivSqrt_io_in_bits_isDiv),
    .io_out_ready(fracDivSqrt_io_out_ready),
    .io_out_valid(fracDivSqrt_io_out_valid),
    .io_out_bits_quot(fracDivSqrt_io_out_bits_quot),
    .io_out_bits_isZeroRem(fracDivSqrt_io_out_bits_isZeroRem)
  );
  RoundingUnit rounding ( // @[FloatDivSqrt.scala 237:24]
    .io_in_rm(rounding_io_in_rm),
    .io_in_frac(rounding_io_in_frac),
    .io_in_sign(rounding_io_in_sign),
    .io_in_guard(rounding_io_in_guard),
    .io_in_round(rounding_io_in_round),
    .io_in_sticky(rounding_io_in_sticky),
    .io_out_fracRounded(rounding_io_out_fracRounded),
    .io_out_fracCout(rounding_io_out_fracCout)
  );
  assign io_in_ready = state == 3'h0; // @[FloatDivSqrt.scala 331:24]
  assign io_out_valid = state == 3'h5; // @[FloatDivSqrt.scala 332:25]
  assign io_out_bits_result = specialCaseReg ? specialResult : commonResult; // @[FloatDivSqrt.scala 333:28]
  assign classify_a_io_in = io_in_bits_a; // @[FloatDivSqrt.scala 120:20]
  assign classify_b_io_in = io_in_bits_b; // @[FloatDivSqrt.scala 123:20]
  assign fracDivSqrt_clock = clock;
  assign fracDivSqrt_reset = reset;
  assign fracDivSqrt_io_in_valid = state == 3'h2; // @[FloatDivSqrt.scala 207:36]
  assign fracDivSqrt_io_in_bits_a = isDivReg | aIsOddExp ? _fracDivSqrt_io_in_bits_a_T_1 : _fracDivSqrt_io_in_bits_a_T_2
    ; // @[FloatDivSqrt.scala 210:34]
  assign fracDivSqrt_io_in_bits_b = {bFracReg,4'h0}; // @[Cat.scala 31:58]
  assign fracDivSqrt_io_in_bits_isDiv = isDivReg; // @[FloatDivSqrt.scala 215:32]
  assign fracDivSqrt_io_out_ready = 1'h1; // @[FloatDivSqrt.scala 206:28]
  assign rounding_io_in_rm = rmReg; // @[FloatDivSqrt.scala 238:21]
  assign rounding_io_in_frac = aFracReg; // @[FloatDivSqrt.scala 239:23]
  assign rounding_io_in_sign = resSignReg; // @[FloatDivSqrt.scala 240:23]
  assign rounding_io_in_guard = gReg; // @[FloatDivSqrt.scala 241:24]
  assign rounding_io_in_round = rReg; // @[FloatDivSqrt.scala 242:24]
  assign rounding_io_in_sticky = sReg; // @[FloatDivSqrt.scala 243:25]
  always @(posedge clock) begin
    if (reset) begin // @[FloatDivSqrt.scala 110:22]
      state <= 3'h0; // @[FloatDivSqrt.scala 110:22]
    end else if (3'h0 == state) begin // @[FloatDivSqrt.scala 275:16]
      if (_rmReg_T) begin // @[FloatDivSqrt.scala 277:25]
        if (sqrtSpecial | divSpecial) begin // @[FloatDivSqrt.scala 278:40]
          state <= 3'h5; // @[FloatDivSqrt.scala 279:17]
        end else begin
          state <= _GEN_16;
        end
      end
    end else if (3'h1 == state) begin // @[FloatDivSqrt.scala 275:16]
      state <= 3'h2; // @[FloatDivSqrt.scala 287:23]
    end else if (3'h2 == state) begin // @[FloatDivSqrt.scala 275:16]
      state <= 3'h3; // @[FloatDivSqrt.scala 288:24]
    end else begin
      state <= _GEN_23;
    end
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      rmReg <= io_in_bits_rm; // @[Reg.scala 17:22]
    end
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      isDivReg <= isDiv; // @[Reg.scala 17:22]
    end
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      resSignReg <= resSign; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[FloatDivSqrt.scala 296:16]
      if (_rmReg_T) begin // @[FloatDivSqrt.scala 298:25]
        aExpReg <= {{1{aExp[8]}},aExp}; // @[FloatDivSqrt.scala 299:17]
      end
    end else if (_T_4) begin // @[FloatDivSqrt.scala 296:16]
      if (aIsSubnormalReg) begin // @[FloatDivSqrt.scala 306:28]
        aExpReg <= _aExpReg_T_3; // @[FloatDivSqrt.scala 307:17]
      end
    end else if (_T_5) begin // @[FloatDivSqrt.scala 296:16]
      if (isDivReg) begin // @[FloatDivSqrt.scala 316:21]
        aExpReg <= _aExpReg_T_6;
      end else begin
        aExpReg <= {{1{_aExpReg_T_10[8]}},_aExpReg_T_10};
      end
    end else if (_T_6) begin // @[FloatDivSqrt.scala 296:16]
      aExpReg <= _GEN_35;
    end else begin
      aExpReg <= _GEN_37;
    end
    aFracReg <= _GEN_48[23:0];
    if (_T) begin // @[FloatDivSqrt.scala 296:16]
      if (_rmReg_T) begin // @[FloatDivSqrt.scala 298:25]
        bExpReg <= {{1{bExp[8]}},bExp}; // @[FloatDivSqrt.scala 301:17]
      end
    end else if (_T_4) begin // @[FloatDivSqrt.scala 296:16]
      if (bIsSubnormalReg) begin // @[FloatDivSqrt.scala 310:28]
        bExpReg <= _bExpReg_T_3; // @[FloatDivSqrt.scala 311:17]
      end
    end
    bFracReg <= _GEN_50[23:0];
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      aIsSubnormalReg <= classify_a_io_isSubnormal; // @[Reg.scala 17:22]
    end
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      bIsSubnormalReg <= classify_b_io_isSubnormal; // @[Reg.scala 17:22]
    end
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      specialCaseReg <= specialCase; // @[Reg.scala 17:22]
    end
    if (_rmReg_T) begin // @[Reg.scala 17:18]
      if (sel_NaN) begin // @[FloatDivSqrt.scala 192:8]
        specialResult <= 32'h7fc00000;
      end else if (sel_Zero) begin // @[FloatDivSqrt.scala 194:10]
        specialResult <= _specialResult_T_3;
      end else begin
        specialResult <= _specialResult_T_7;
      end
    end
    gReg <= fracShifted[2]; // @[FloatDivSqrt.scala 229:46]
    rReg <= fracShifted[1]; // @[FloatDivSqrt.scala 230:48]
    sReg <= ~fracDivSqrt_io_out_bits_isZeroRem | |fracShifted[0]; // @[FloatDivSqrt.scala 231:46]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  rmReg = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  isDivReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  resSignReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  aExpReg = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  aFracReg = _RAND_5[23:0];
  _RAND_6 = {1{`RANDOM}};
  bExpReg = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  bFracReg = _RAND_7[23:0];
  _RAND_8 = {1{`RANDOM}};
  aIsSubnormalReg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  bIsSubnormalReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  specialCaseReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  specialResult = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  gReg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rReg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sReg = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_9(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits = io_in_0_valid ? io_in_0_bits : io_in_1_bits; // @[Arbiter.scala 139:15 141:26 143:19]
endmodule
module SFUexe(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_in1_0,
  input  [31:0] io_in_bits_in1_1,
  input  [31:0] io_in_bits_in1_2,
  input  [31:0] io_in_bits_in1_3,
  input  [31:0] io_in_bits_in1_4,
  input  [31:0] io_in_bits_in1_5,
  input  [31:0] io_in_bits_in1_6,
  input  [31:0] io_in_bits_in1_7,
  input  [31:0] io_in_bits_in2_0,
  input  [31:0] io_in_bits_in2_1,
  input  [31:0] io_in_bits_in2_2,
  input  [31:0] io_in_bits_in2_3,
  input  [31:0] io_in_bits_in2_4,
  input  [31:0] io_in_bits_in2_5,
  input  [31:0] io_in_bits_in2_6,
  input  [31:0] io_in_bits_in2_7,
  input         io_in_bits_mask_0,
  input         io_in_bits_mask_1,
  input         io_in_bits_mask_2,
  input         io_in_bits_mask_3,
  input         io_in_bits_mask_4,
  input         io_in_bits_mask_5,
  input         io_in_bits_mask_6,
  input         io_in_bits_mask_7,
  input  [1:0]  io_in_bits_ctrl_wid,
  input         io_in_bits_ctrl_fp,
  input         io_in_bits_ctrl_reverse,
  input         io_in_bits_ctrl_isvec,
  input  [5:0]  io_in_bits_ctrl_alu_fn,
  input  [4:0]  io_in_bits_ctrl_reg_idxw,
  input         io_in_bits_ctrl_wfd,
  input         io_in_bits_ctrl_wxd,
  input  [2:0]  io_rm,
  input         io_out_x_ready,
  output        io_out_x_valid,
  output [31:0] io_out_x_bits_wb_wxd_rd,
  output        io_out_x_bits_wxd,
  output [4:0]  io_out_x_bits_reg_idxw,
  output [1:0]  io_out_x_bits_warp_id,
  input         io_out_v_ready,
  output        io_out_v_valid,
  output [31:0] io_out_v_bits_wb_wfd_rd_0,
  output [31:0] io_out_v_bits_wb_wfd_rd_1,
  output [31:0] io_out_v_bits_wb_wfd_rd_2,
  output [31:0] io_out_v_bits_wb_wfd_rd_3,
  output [31:0] io_out_v_bits_wb_wfd_rd_4,
  output [31:0] io_out_v_bits_wb_wfd_rd_5,
  output [31:0] io_out_v_bits_wb_wfd_rd_6,
  output [31:0] io_out_v_bits_wb_wfd_rd_7,
  output        io_out_v_bits_wfd_mask_0,
  output        io_out_v_bits_wfd_mask_1,
  output        io_out_v_bits_wfd_mask_2,
  output        io_out_v_bits_wfd_mask_3,
  output        io_out_v_bits_wfd_mask_4,
  output        io_out_v_bits_wfd_mask_5,
  output        io_out_v_bits_wfd_mask_6,
  output        io_out_v_bits_wfd_mask_7,
  output        io_out_v_bits_wfd,
  output [4:0]  io_out_v_bits_reg_idxw,
  output [1:0]  io_out_v_bits_warp_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  result_x_clock; // @[execution.scala 176:22]
  wire  result_x_reset; // @[execution.scala 176:22]
  wire  result_x_io_enq_ready; // @[execution.scala 176:22]
  wire  result_x_io_enq_valid; // @[execution.scala 176:22]
  wire [31:0] result_x_io_enq_bits_wb_wxd_rd; // @[execution.scala 176:22]
  wire  result_x_io_enq_bits_wxd; // @[execution.scala 176:22]
  wire [4:0] result_x_io_enq_bits_reg_idxw; // @[execution.scala 176:22]
  wire [1:0] result_x_io_enq_bits_warp_id; // @[execution.scala 176:22]
  wire  result_x_io_deq_ready; // @[execution.scala 176:22]
  wire  result_x_io_deq_valid; // @[execution.scala 176:22]
  wire [31:0] result_x_io_deq_bits_wb_wxd_rd; // @[execution.scala 176:22]
  wire  result_x_io_deq_bits_wxd; // @[execution.scala 176:22]
  wire [4:0] result_x_io_deq_bits_reg_idxw; // @[execution.scala 176:22]
  wire [1:0] result_x_io_deq_bits_warp_id; // @[execution.scala 176:22]
  wire  result_v_clock; // @[execution.scala 177:22]
  wire  result_v_reset; // @[execution.scala 177:22]
  wire  result_v_io_enq_ready; // @[execution.scala 177:22]
  wire  result_v_io_enq_valid; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_0; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_1; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_2; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_3; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_4; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_5; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_6; // @[execution.scala 177:22]
  wire [31:0] result_v_io_enq_bits_wb_wfd_rd_7; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_0; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_1; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_2; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_3; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_4; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_5; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_6; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd_mask_7; // @[execution.scala 177:22]
  wire  result_v_io_enq_bits_wfd; // @[execution.scala 177:22]
  wire [4:0] result_v_io_enq_bits_reg_idxw; // @[execution.scala 177:22]
  wire [1:0] result_v_io_enq_bits_warp_id; // @[execution.scala 177:22]
  wire  result_v_io_deq_ready; // @[execution.scala 177:22]
  wire  result_v_io_deq_valid; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_0; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_1; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_2; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_3; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_4; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_5; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_6; // @[execution.scala 177:22]
  wire [31:0] result_v_io_deq_bits_wb_wfd_rd_7; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_0; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_1; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_2; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_3; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_4; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_5; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_6; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd_mask_7; // @[execution.scala 177:22]
  wire  result_v_io_deq_bits_wfd; // @[execution.scala 177:22]
  wire [4:0] result_v_io_deq_bits_reg_idxw; // @[execution.scala 177:22]
  wire [1:0] result_v_io_deq_bits_warp_id; // @[execution.scala 177:22]
  wire  data_buffer_clock; // @[Decoupled.scala 361:21]
  wire  data_buffer_reset; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_0; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_1; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_2; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_3; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_4; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_5; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_6; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in1_7; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_0; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_1; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_2; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_3; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_4; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_5; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_6; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_enq_bits_in2_7; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_0; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_1; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_2; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_3; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_4; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_5; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_6; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_mask_7; // @[Decoupled.scala 361:21]
  wire [1:0] data_buffer_io_enq_bits_ctrl_wid; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_ctrl_fp; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_ctrl_reverse; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_ctrl_isvec; // @[Decoupled.scala 361:21]
  wire [5:0] data_buffer_io_enq_bits_ctrl_alu_fn; // @[Decoupled.scala 361:21]
  wire [4:0] data_buffer_io_enq_bits_ctrl_reg_idxw; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_ctrl_wfd; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_enq_bits_ctrl_wxd; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_0; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_1; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_2; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_3; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_4; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_5; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_6; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in1_7; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_0; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_1; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_2; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_3; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_4; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_5; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_6; // @[Decoupled.scala 361:21]
  wire [31:0] data_buffer_io_deq_bits_in2_7; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_0; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_1; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_2; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_3; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_4; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_5; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_6; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_mask_7; // @[Decoupled.scala 361:21]
  wire [1:0] data_buffer_io_deq_bits_ctrl_wid; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_ctrl_fp; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_ctrl_reverse; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_ctrl_isvec; // @[Decoupled.scala 361:21]
  wire [5:0] data_buffer_io_deq_bits_ctrl_alu_fn; // @[Decoupled.scala 361:21]
  wire [4:0] data_buffer_io_deq_bits_ctrl_reg_idxw; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_ctrl_wfd; // @[Decoupled.scala 361:21]
  wire  data_buffer_io_deq_bits_ctrl_wxd; // @[Decoupled.scala 361:21]
  wire  IntDivMod_clock; // @[execution.scala 209:46]
  wire  IntDivMod_reset; // @[execution.scala 209:46]
  wire  IntDivMod_io_in_ready; // @[execution.scala 209:46]
  wire  IntDivMod_io_in_valid; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_io_in_bits_a; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_io_in_bits_d; // @[execution.scala 209:46]
  wire  IntDivMod_io_in_bits_signed; // @[execution.scala 209:46]
  wire  IntDivMod_io_out_ready; // @[execution.scala 209:46]
  wire  IntDivMod_io_out_valid; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_io_out_bits_q; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_io_out_bits_r; // @[execution.scala 209:46]
  wire  IntDivMod_1_clock; // @[execution.scala 209:46]
  wire  IntDivMod_1_reset; // @[execution.scala 209:46]
  wire  IntDivMod_1_io_in_ready; // @[execution.scala 209:46]
  wire  IntDivMod_1_io_in_valid; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_1_io_in_bits_a; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_1_io_in_bits_d; // @[execution.scala 209:46]
  wire  IntDivMod_1_io_in_bits_signed; // @[execution.scala 209:46]
  wire  IntDivMod_1_io_out_ready; // @[execution.scala 209:46]
  wire  IntDivMod_1_io_out_valid; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_1_io_out_bits_q; // @[execution.scala 209:46]
  wire [31:0] IntDivMod_1_io_out_bits_r; // @[execution.scala 209:46]
  wire  FloatDivSqrt_clock; // @[execution.scala 210:48]
  wire  FloatDivSqrt_reset; // @[execution.scala 210:48]
  wire  FloatDivSqrt_io_in_ready; // @[execution.scala 210:48]
  wire  FloatDivSqrt_io_in_valid; // @[execution.scala 210:48]
  wire [2:0] FloatDivSqrt_io_in_bits_op; // @[execution.scala 210:48]
  wire [31:0] FloatDivSqrt_io_in_bits_a; // @[execution.scala 210:48]
  wire [31:0] FloatDivSqrt_io_in_bits_b; // @[execution.scala 210:48]
  wire [2:0] FloatDivSqrt_io_in_bits_rm; // @[execution.scala 210:48]
  wire  FloatDivSqrt_io_out_ready; // @[execution.scala 210:48]
  wire  FloatDivSqrt_io_out_valid; // @[execution.scala 210:48]
  wire [31:0] FloatDivSqrt_io_out_bits_result; // @[execution.scala 210:48]
  wire  FloatDivSqrt_1_clock; // @[execution.scala 210:48]
  wire  FloatDivSqrt_1_reset; // @[execution.scala 210:48]
  wire  FloatDivSqrt_1_io_in_ready; // @[execution.scala 210:48]
  wire  FloatDivSqrt_1_io_in_valid; // @[execution.scala 210:48]
  wire [2:0] FloatDivSqrt_1_io_in_bits_op; // @[execution.scala 210:48]
  wire [31:0] FloatDivSqrt_1_io_in_bits_a; // @[execution.scala 210:48]
  wire [31:0] FloatDivSqrt_1_io_in_bits_b; // @[execution.scala 210:48]
  wire [2:0] FloatDivSqrt_1_io_in_bits_rm; // @[execution.scala 210:48]
  wire  FloatDivSqrt_1_io_out_ready; // @[execution.scala 210:48]
  wire  FloatDivSqrt_1_io_out_valid; // @[execution.scala 210:48]
  wire [31:0] FloatDivSqrt_1_io_out_bits_result; // @[execution.scala 210:48]
  wire  Arbiter_io_in_0_ready; // @[execution.scala 211:55]
  wire  Arbiter_io_in_0_valid; // @[execution.scala 211:55]
  wire [31:0] Arbiter_io_in_0_bits; // @[execution.scala 211:55]
  wire  Arbiter_io_in_1_ready; // @[execution.scala 211:55]
  wire  Arbiter_io_in_1_valid; // @[execution.scala 211:55]
  wire [31:0] Arbiter_io_in_1_bits; // @[execution.scala 211:55]
  wire  Arbiter_io_out_ready; // @[execution.scala 211:55]
  wire  Arbiter_io_out_valid; // @[execution.scala 211:55]
  wire [31:0] Arbiter_io_out_bits; // @[execution.scala 211:55]
  wire  Arbiter_1_io_in_0_ready; // @[execution.scala 211:55]
  wire  Arbiter_1_io_in_0_valid; // @[execution.scala 211:55]
  wire [31:0] Arbiter_1_io_in_0_bits; // @[execution.scala 211:55]
  wire  Arbiter_1_io_in_1_ready; // @[execution.scala 211:55]
  wire  Arbiter_1_io_in_1_valid; // @[execution.scala 211:55]
  wire [31:0] Arbiter_1_io_in_1_bits; // @[execution.scala 211:55]
  wire  Arbiter_1_io_out_ready; // @[execution.scala 211:55]
  wire  Arbiter_1_io_out_valid; // @[execution.scala 211:55]
  wire [31:0] Arbiter_1_io_out_bits; // @[execution.scala 211:55]
  reg [1:0] state; // @[execution.scala 179:20]
  reg [7:0] mask; // @[execution.scala 182:19]
  wire  mask_grp_0 = |mask[1:0]; // @[execution.scala 185:86]
  wire  mask_grp_1 = |mask[3:2]; // @[execution.scala 185:86]
  wire  mask_grp_2 = |mask[5:4]; // @[execution.scala 185:86]
  reg [31:0] out_data_0; // @[execution.scala 189:23]
  reg [31:0] out_data_1; // @[execution.scala 189:23]
  reg [31:0] out_data_2; // @[execution.scala 189:23]
  reg [31:0] out_data_3; // @[execution.scala 189:23]
  reg [31:0] out_data_4; // @[execution.scala 189:23]
  reg [31:0] out_data_5; // @[execution.scala 189:23]
  reg [31:0] out_data_6; // @[execution.scala 189:23]
  reg [31:0] out_data_7; // @[execution.scala 189:23]
  wire [1:0] _i_cnt_T = mask_grp_2 ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _i_cnt_T_1 = mask_grp_1 ? 2'h1 : _i_cnt_T; // @[Mux.scala 47:70]
  wire [1:0] i_cnt = mask_grp_0 ? 2'h0 : _i_cnt_T_1; // @[Mux.scala 47:70]
  reg  i_valid; // @[execution.scala 193:24]
  wire  _T = 2'h0 == i_cnt; // @[execution.scala 200:18]
  wire [31:0] i_2__0 = data_buffer_io_deq_bits_in2_0; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1__0 = data_buffer_io_deq_bits_in1_0; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_1_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_2__0 : i_1__0; // @[execution.scala 203:19]
  wire [31:0] i_2__1 = data_buffer_io_deq_bits_in2_1; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1__1 = data_buffer_io_deq_bits_in1_1; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_1_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_2__1 : i_1__1; // @[execution.scala 203:19]
  wire [31:0] _T_2_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_1__0 : i_2__0; // @[execution.scala 204:19]
  wire [31:0] _T_2_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_1__1 : i_2__1; // @[execution.scala 204:19]
  wire [31:0] _GEN_0 = 2'h0 == i_cnt ? _T_1_0 : 32'h0; // @[execution.scala 200:27 203:14]
  wire [31:0] _GEN_1 = 2'h0 == i_cnt ? _T_1_1 : 32'h0; // @[execution.scala 200:27 203:14]
  wire [31:0] _GEN_2 = 2'h0 == i_cnt ? _T_2_0 : 32'h0; // @[execution.scala 200:27 204:14]
  wire [31:0] _GEN_3 = 2'h0 == i_cnt ? _T_2_1 : 32'h0; // @[execution.scala 200:27 204:14]
  wire  _T_6 = 2'h1 == i_cnt; // @[execution.scala 200:18]
  wire [31:0] i_2_1_0 = data_buffer_io_deq_bits_in2_2; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1_1_0 = data_buffer_io_deq_bits_in1_2; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_7_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_2_1_0 : i_1_1_0; // @[execution.scala 203:19]
  wire [31:0] i_2_1_1 = data_buffer_io_deq_bits_in2_3; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1_1_1 = data_buffer_io_deq_bits_in1_3; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_7_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_2_1_1 : i_1_1_1; // @[execution.scala 203:19]
  wire [31:0] _T_8_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_1_1_0 : i_2_1_0; // @[execution.scala 204:19]
  wire [31:0] _T_8_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_1_1_1 : i_2_1_1; // @[execution.scala 204:19]
  wire [31:0] _GEN_8 = 2'h1 == i_cnt ? _T_7_0 : _GEN_0; // @[execution.scala 200:27 203:14]
  wire [31:0] _GEN_9 = 2'h1 == i_cnt ? _T_7_1 : _GEN_1; // @[execution.scala 200:27 203:14]
  wire [31:0] _GEN_10 = 2'h1 == i_cnt ? _T_8_0 : _GEN_2; // @[execution.scala 200:27 204:14]
  wire [31:0] _GEN_11 = 2'h1 == i_cnt ? _T_8_1 : _GEN_3; // @[execution.scala 200:27 204:14]
  wire  _GEN_14 = 2'h1 == i_cnt ? mask[2] : 2'h0 == i_cnt & mask[0]; // @[execution.scala 200:27 206:13]
  wire  _GEN_15 = 2'h1 == i_cnt ? mask[3] : 2'h0 == i_cnt & mask[1]; // @[execution.scala 200:27 206:13]
  wire  _T_12 = 2'h2 == i_cnt; // @[execution.scala 200:18]
  wire [31:0] i_2_2_0 = data_buffer_io_deq_bits_in2_4; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1_2_0 = data_buffer_io_deq_bits_in1_4; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_13_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_2_2_0 : i_1_2_0; // @[execution.scala 203:19]
  wire [31:0] i_2_2_1 = data_buffer_io_deq_bits_in2_5; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1_2_1 = data_buffer_io_deq_bits_in1_5; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_13_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_2_2_1 : i_1_2_1; // @[execution.scala 203:19]
  wire [31:0] _T_14_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_1_2_0 : i_2_2_0; // @[execution.scala 204:19]
  wire [31:0] _T_14_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_1_2_1 : i_2_2_1; // @[execution.scala 204:19]
  wire [31:0] _GEN_16 = 2'h2 == i_cnt ? _T_13_0 : _GEN_8; // @[execution.scala 200:27 203:14]
  wire [31:0] _GEN_17 = 2'h2 == i_cnt ? _T_13_1 : _GEN_9; // @[execution.scala 200:27 203:14]
  wire [31:0] _GEN_18 = 2'h2 == i_cnt ? _T_14_0 : _GEN_10; // @[execution.scala 200:27 204:14]
  wire [31:0] _GEN_19 = 2'h2 == i_cnt ? _T_14_1 : _GEN_11; // @[execution.scala 200:27 204:14]
  wire  _GEN_22 = 2'h2 == i_cnt ? mask[4] : _GEN_14; // @[execution.scala 200:27 206:13]
  wire  _GEN_23 = 2'h2 == i_cnt ? mask[5] : _GEN_15; // @[execution.scala 200:27 206:13]
  wire  _T_18 = 2'h3 == i_cnt; // @[execution.scala 200:18]
  wire [31:0] i_2_3_0 = data_buffer_io_deq_bits_in2_6; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1_3_0 = data_buffer_io_deq_bits_in1_6; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_19_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_2_3_0 : i_1_3_0; // @[execution.scala 203:19]
  wire [31:0] i_2_3_1 = data_buffer_io_deq_bits_in2_7; // @[execution.scala 202:{24,24}]
  wire [31:0] i_1_3_1 = data_buffer_io_deq_bits_in1_7; // @[execution.scala 201:{24,24}]
  wire [31:0] _T_19_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_2_3_1 : i_1_3_1; // @[execution.scala 203:19]
  wire [31:0] _T_20_0 = data_buffer_io_deq_bits_ctrl_reverse ? i_1_3_0 : i_2_3_0; // @[execution.scala 204:19]
  wire [31:0] _T_20_1 = data_buffer_io_deq_bits_ctrl_reverse ? i_1_3_1 : i_2_3_1; // @[execution.scala 204:19]
  wire [31:0] i_data1_0 = 2'h3 == i_cnt ? _T_19_0 : _GEN_16; // @[execution.scala 200:27 203:14]
  wire [31:0] i_data1_1 = 2'h3 == i_cnt ? _T_19_1 : _GEN_17; // @[execution.scala 200:27 203:14]
  wire [31:0] i_data2_0 = 2'h3 == i_cnt ? _T_20_0 : _GEN_18; // @[execution.scala 200:27 204:14]
  wire [31:0] i_data2_1 = 2'h3 == i_cnt ? _T_20_1 : _GEN_19; // @[execution.scala 200:27 204:14]
  wire  i_mask_0 = 2'h3 == i_cnt ? mask[6] : _GEN_22; // @[execution.scala 200:27 206:13]
  wire  i_mask_1 = 2'h3 == i_cnt ? mask[7] : _GEN_23; // @[execution.scala 200:27 206:13]
  wire  alu_out_arbiter_0_out_valid = Arbiter_io_out_valid; // @[execution.scala 211:{30,30}]
  wire  alu_out_arbiter_1_out_valid = Arbiter_1_io_out_valid; // @[execution.scala 211:{30,30}]
  wire  alu_out_arbiter_0_out_ready = alu_out_arbiter_0_out_valid & alu_out_arbiter_1_out_valid; // @[execution.scala 212:87]
  wire  _result_x_io_enq_valid_T = state == 2'h2; // @[execution.scala 225:31]
  wire  o_ready = data_buffer_io_deq_bits_ctrl_isvec & result_v_io_enq_ready | ~data_buffer_io_deq_bits_ctrl_isvec &
    result_x_io_enq_ready; // @[execution.scala 227:51]
  wire [31:0] intDiv_0_out_bits_r = IntDivMod_io_out_bits_r; // @[execution.scala 209:{21,21}]
  wire [31:0] intDiv_0_out_bits_q = IntDivMod_io_out_bits_q; // @[execution.scala 209:{21,21}]
  wire [31:0] _GEN_32 = _T & i_mask_0 ? i_data1_0 : 32'h1; // @[execution.scala 237:25 243:41 244:25]
  wire [31:0] _GEN_33 = _T & i_mask_0 ? i_data2_0 : 32'h1; // @[execution.scala 238:25 243:41 245:25]
  wire [31:0] _GEN_34 = _T & i_mask_0 ? i_data1_0 : 32'h3f800000; // @[execution.scala 239:27 243:41 246:27]
  wire [31:0] _GEN_35 = _T & i_mask_0 ? i_data2_0 : 32'h3f800000; // @[execution.scala 240:27 243:41 247:27]
  wire [31:0] _GEN_37 = _T_6 & i_mask_0 ? i_data1_0 : _GEN_32; // @[execution.scala 243:41 244:25]
  wire [31:0] _GEN_38 = _T_6 & i_mask_0 ? i_data2_0 : _GEN_33; // @[execution.scala 243:41 245:25]
  wire [31:0] _GEN_39 = _T_6 & i_mask_0 ? i_data1_0 : _GEN_34; // @[execution.scala 243:41 246:27]
  wire [31:0] _GEN_40 = _T_6 & i_mask_0 ? i_data2_0 : _GEN_35; // @[execution.scala 243:41 247:27]
  wire [31:0] _GEN_42 = _T_12 & i_mask_0 ? i_data1_0 : _GEN_37; // @[execution.scala 243:41 244:25]
  wire [31:0] _GEN_43 = _T_12 & i_mask_0 ? i_data2_0 : _GEN_38; // @[execution.scala 243:41 245:25]
  wire [31:0] _GEN_44 = _T_12 & i_mask_0 ? i_data1_0 : _GEN_39; // @[execution.scala 243:41 246:27]
  wire [31:0] _GEN_45 = _T_12 & i_mask_0 ? i_data2_0 : _GEN_40; // @[execution.scala 243:41 247:27]
  wire [31:0] intDiv_1_out_bits_r = IntDivMod_1_io_out_bits_r; // @[execution.scala 209:{21,21}]
  wire [31:0] intDiv_1_out_bits_q = IntDivMod_1_io_out_bits_q; // @[execution.scala 209:{21,21}]
  wire [31:0] _GEN_52 = _T & i_mask_1 ? i_data1_1 : 32'h1; // @[execution.scala 237:25 243:41 244:25]
  wire [31:0] _GEN_53 = _T & i_mask_1 ? i_data2_1 : 32'h1; // @[execution.scala 238:25 243:41 245:25]
  wire [31:0] _GEN_54 = _T & i_mask_1 ? i_data1_1 : 32'h3f800000; // @[execution.scala 239:27 243:41 246:27]
  wire [31:0] _GEN_55 = _T & i_mask_1 ? i_data2_1 : 32'h3f800000; // @[execution.scala 240:27 243:41 247:27]
  wire [31:0] _GEN_57 = _T_6 & i_mask_1 ? i_data1_1 : _GEN_52; // @[execution.scala 243:41 244:25]
  wire [31:0] _GEN_58 = _T_6 & i_mask_1 ? i_data2_1 : _GEN_53; // @[execution.scala 243:41 245:25]
  wire [31:0] _GEN_59 = _T_6 & i_mask_1 ? i_data1_1 : _GEN_54; // @[execution.scala 243:41 246:27]
  wire [31:0] _GEN_60 = _T_6 & i_mask_1 ? i_data2_1 : _GEN_55; // @[execution.scala 243:41 247:27]
  wire [31:0] _GEN_62 = _T_12 & i_mask_1 ? i_data1_1 : _GEN_57; // @[execution.scala 243:41 244:25]
  wire [31:0] _GEN_63 = _T_12 & i_mask_1 ? i_data2_1 : _GEN_58; // @[execution.scala 243:41 245:25]
  wire [31:0] _GEN_64 = _T_12 & i_mask_1 ? i_data1_1 : _GEN_59; // @[execution.scala 243:41 246:27]
  wire [31:0] _GEN_65 = _T_12 & i_mask_1 ? i_data2_1 : _GEN_60; // @[execution.scala 243:41 247:27]
  wire  floatDiv_0_in_ready = FloatDivSqrt_io_in_ready; // @[execution.scala 210:{23,23}]
  wire  intDiv_0_in_ready = IntDivMod_io_in_ready; // @[execution.scala 209:{21,21}]
  wire  i_ready = data_buffer_io_deq_bits_ctrl_fp ? floatDiv_0_in_ready : intDiv_0_in_ready; // @[execution.scala 256:22]
  wire  alu_out_fire = alu_out_arbiter_0_out_ready & alu_out_arbiter_0_out_valid; // @[Decoupled.scala 50:35]
  wire  _T_41 = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  wire [7:0] _mask_T = {io_in_bits_mask_7,io_in_bits_mask_6,io_in_bits_mask_5,io_in_bits_mask_4,io_in_bits_mask_3,
    io_in_bits_mask_2,io_in_bits_mask_1,io_in_bits_mask_0}; // @[execution.scala 264:31]
  wire [7:0] _GEN_73 = _T_41 ? _mask_T : mask; // @[execution.scala 262:25 264:13 182:19]
  wire  _GEN_74 = _T_41 | i_valid; // @[execution.scala 262:25 265:16 193:24]
  wire  _GEN_75 = i_valid & i_ready ? 1'h0 : i_valid; // @[execution.scala 269:30 270:16 193:24]
  wire [31:0] _GEN_159 = {{24'd0}, mask}; // @[execution.scala 275:32]
  wire [31:0] next_mask = _GEN_159 & 32'hfffffffc; // @[execution.scala 275:32]
  wire [1:0] _GEN_76 = ~(|next_mask) ? 2'h2 : state; // @[execution.scala 179:20 279:35 280:21]
  wire  _GEN_77 = ~(|next_mask) ? 1'h0 : 1'h1; // @[execution.scala 277:20 279:35 281:22]
  wire [31:0] _GEN_78 = _T ? next_mask : {{24'd0}, mask}; // @[execution.scala 274:33 276:18 182:19]
  wire  _GEN_79 = _T ? _GEN_77 : _GEN_75; // @[execution.scala 274:33]
  wire [31:0] alu_out_arbiter_0_out_bits = Arbiter_io_out_bits; // @[execution.scala 211:{30,30}]
  wire [31:0] _GEN_80 = _T ? alu_out_arbiter_0_out_bits : out_data_0; // @[execution.scala 189:23 274:33 278:61]
  wire [31:0] alu_out_arbiter_1_out_bits = Arbiter_1_io_out_bits; // @[execution.scala 211:{30,30}]
  wire [31:0] _GEN_81 = _T ? alu_out_arbiter_1_out_bits : out_data_1; // @[execution.scala 189:23 274:33 278:61]
  wire [1:0] _GEN_82 = _T ? _GEN_76 : state; // @[execution.scala 179:20 274:33]
  wire [33:0] _GEN_160 = {{26'd0}, mask}; // @[execution.scala 275:32]
  wire [33:0] next_mask_1 = _GEN_160 & 34'h3fffffff3; // @[execution.scala 275:32]
  wire [1:0] _GEN_83 = ~(|next_mask_1) ? 2'h2 : _GEN_82; // @[execution.scala 279:35 280:21]
  wire  _GEN_84 = ~(|next_mask_1) ? 1'h0 : 1'h1; // @[execution.scala 277:20 279:35 281:22]
  wire [33:0] _GEN_85 = _T_6 ? next_mask_1 : {{2'd0}, _GEN_78}; // @[execution.scala 274:33 276:18]
  wire  _GEN_86 = _T_6 ? _GEN_84 : _GEN_79; // @[execution.scala 274:33]
  wire [31:0] _GEN_87 = _T_6 ? alu_out_arbiter_0_out_bits : out_data_2; // @[execution.scala 189:23 274:33 278:61]
  wire [31:0] _GEN_88 = _T_6 ? alu_out_arbiter_1_out_bits : out_data_3; // @[execution.scala 189:23 274:33 278:61]
  wire [1:0] _GEN_89 = _T_6 ? _GEN_83 : _GEN_82; // @[execution.scala 274:33]
  wire [35:0] _GEN_161 = {{28'd0}, mask}; // @[execution.scala 275:32]
  wire [35:0] next_mask_2 = _GEN_161 & 36'hfffffffcf; // @[execution.scala 275:32]
  wire [1:0] _GEN_90 = ~(|next_mask_2) ? 2'h2 : _GEN_89; // @[execution.scala 279:35 280:21]
  wire  _GEN_91 = ~(|next_mask_2) ? 1'h0 : 1'h1; // @[execution.scala 277:20 279:35 281:22]
  wire [35:0] _GEN_92 = _T_12 ? next_mask_2 : {{2'd0}, _GEN_85}; // @[execution.scala 274:33 276:18]
  wire  _GEN_93 = _T_12 ? _GEN_91 : _GEN_86; // @[execution.scala 274:33]
  wire [31:0] _GEN_94 = _T_12 ? alu_out_arbiter_0_out_bits : out_data_4; // @[execution.scala 189:23 274:33 278:61]
  wire [31:0] _GEN_95 = _T_12 ? alu_out_arbiter_1_out_bits : out_data_5; // @[execution.scala 189:23 274:33 278:61]
  wire [1:0] _GEN_96 = _T_12 ? _GEN_90 : _GEN_89; // @[execution.scala 274:33]
  wire [37:0] _GEN_162 = {{30'd0}, mask}; // @[execution.scala 275:32]
  wire [37:0] next_mask_3 = _GEN_162 & 38'h3fffffff3f; // @[execution.scala 275:32]
  wire [1:0] _GEN_97 = ~(|next_mask_3) ? 2'h2 : _GEN_96; // @[execution.scala 279:35 280:21]
  wire  _GEN_98 = ~(|next_mask_3) ? 1'h0 : 1'h1; // @[execution.scala 277:20 279:35 281:22]
  wire [37:0] _GEN_99 = _T_18 ? next_mask_3 : {{2'd0}, _GEN_92}; // @[execution.scala 274:33 276:18]
  wire  _GEN_100 = _T_18 ? _GEN_98 : _GEN_93; // @[execution.scala 274:33]
  wire [31:0] _GEN_101 = _T_18 ? alu_out_arbiter_0_out_bits : out_data_6; // @[execution.scala 189:23 274:33 278:61]
  wire [31:0] _GEN_102 = _T_18 ? alu_out_arbiter_1_out_bits : out_data_7; // @[execution.scala 189:23 274:33 278:61]
  wire [1:0] _GEN_103 = _T_18 ? _GEN_97 : _GEN_96; // @[execution.scala 274:33]
  wire [31:0] _GEN_104 = alu_out_fire ? alu_out_arbiter_0_out_bits : out_data_0; // @[execution.scala 287:32 288:21 189:23]
  wire [1:0] _GEN_105 = alu_out_fire ? 2'h2 : state; // @[execution.scala 287:32 289:15 179:20]
  wire  _GEN_106 = alu_out_fire ? 1'h0 : _GEN_75; // @[execution.scala 287:32 290:16]
  wire [37:0] _GEN_107 = data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire ? _GEN_99 : {{30'd0}, mask}; // @[execution.scala 182:19 272:56]
  wire [1:0] _GEN_118 = o_ready ? 2'h0 : state; // @[execution.scala 295:20 296:14 179:20]
  wire [31:0] _GEN_119 = o_ready ? 32'h0 : out_data_0; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_120 = o_ready ? 32'h0 : out_data_1; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_121 = o_ready ? 32'h0 : out_data_2; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_122 = o_ready ? 32'h0 : out_data_3; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_123 = o_ready ? 32'h0 : out_data_4; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_124 = o_ready ? 32'h0 : out_data_5; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_125 = o_ready ? 32'h0 : out_data_6; // @[execution.scala 295:20 297:17 189:23]
  wire [31:0] _GEN_126 = o_ready ? 32'h0 : out_data_7; // @[execution.scala 295:20 297:17 189:23]
  wire [37:0] _GEN_137 = 2'h1 == state ? _GEN_107 : {{30'd0}, mask}; // @[execution.scala 260:16 182:19]
  wire [37:0] _GEN_148 = 2'h0 == state ? {{30'd0}, _GEN_73} : _GEN_137; // @[execution.scala 260:16]
  wire [37:0] _GEN_163 = reset ? 38'h0 : _GEN_148; // @[execution.scala 182:{19,19}]
  Queue_1 result_x ( // @[execution.scala 176:22]
    .clock(result_x_clock),
    .reset(result_x_reset),
    .io_enq_ready(result_x_io_enq_ready),
    .io_enq_valid(result_x_io_enq_valid),
    .io_enq_bits_wb_wxd_rd(result_x_io_enq_bits_wb_wxd_rd),
    .io_enq_bits_wxd(result_x_io_enq_bits_wxd),
    .io_enq_bits_reg_idxw(result_x_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_x_io_enq_bits_warp_id),
    .io_deq_ready(result_x_io_deq_ready),
    .io_deq_valid(result_x_io_deq_valid),
    .io_deq_bits_wb_wxd_rd(result_x_io_deq_bits_wb_wxd_rd),
    .io_deq_bits_wxd(result_x_io_deq_bits_wxd),
    .io_deq_bits_reg_idxw(result_x_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_x_io_deq_bits_warp_id)
  );
  Queue_3 result_v ( // @[execution.scala 177:22]
    .clock(result_v_clock),
    .reset(result_v_reset),
    .io_enq_ready(result_v_io_enq_ready),
    .io_enq_valid(result_v_io_enq_valid),
    .io_enq_bits_wb_wfd_rd_0(result_v_io_enq_bits_wb_wfd_rd_0),
    .io_enq_bits_wb_wfd_rd_1(result_v_io_enq_bits_wb_wfd_rd_1),
    .io_enq_bits_wb_wfd_rd_2(result_v_io_enq_bits_wb_wfd_rd_2),
    .io_enq_bits_wb_wfd_rd_3(result_v_io_enq_bits_wb_wfd_rd_3),
    .io_enq_bits_wb_wfd_rd_4(result_v_io_enq_bits_wb_wfd_rd_4),
    .io_enq_bits_wb_wfd_rd_5(result_v_io_enq_bits_wb_wfd_rd_5),
    .io_enq_bits_wb_wfd_rd_6(result_v_io_enq_bits_wb_wfd_rd_6),
    .io_enq_bits_wb_wfd_rd_7(result_v_io_enq_bits_wb_wfd_rd_7),
    .io_enq_bits_wfd_mask_0(result_v_io_enq_bits_wfd_mask_0),
    .io_enq_bits_wfd_mask_1(result_v_io_enq_bits_wfd_mask_1),
    .io_enq_bits_wfd_mask_2(result_v_io_enq_bits_wfd_mask_2),
    .io_enq_bits_wfd_mask_3(result_v_io_enq_bits_wfd_mask_3),
    .io_enq_bits_wfd_mask_4(result_v_io_enq_bits_wfd_mask_4),
    .io_enq_bits_wfd_mask_5(result_v_io_enq_bits_wfd_mask_5),
    .io_enq_bits_wfd_mask_6(result_v_io_enq_bits_wfd_mask_6),
    .io_enq_bits_wfd_mask_7(result_v_io_enq_bits_wfd_mask_7),
    .io_enq_bits_wfd(result_v_io_enq_bits_wfd),
    .io_enq_bits_reg_idxw(result_v_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_v_io_enq_bits_warp_id),
    .io_deq_ready(result_v_io_deq_ready),
    .io_deq_valid(result_v_io_deq_valid),
    .io_deq_bits_wb_wfd_rd_0(result_v_io_deq_bits_wb_wfd_rd_0),
    .io_deq_bits_wb_wfd_rd_1(result_v_io_deq_bits_wb_wfd_rd_1),
    .io_deq_bits_wb_wfd_rd_2(result_v_io_deq_bits_wb_wfd_rd_2),
    .io_deq_bits_wb_wfd_rd_3(result_v_io_deq_bits_wb_wfd_rd_3),
    .io_deq_bits_wb_wfd_rd_4(result_v_io_deq_bits_wb_wfd_rd_4),
    .io_deq_bits_wb_wfd_rd_5(result_v_io_deq_bits_wb_wfd_rd_5),
    .io_deq_bits_wb_wfd_rd_6(result_v_io_deq_bits_wb_wfd_rd_6),
    .io_deq_bits_wb_wfd_rd_7(result_v_io_deq_bits_wb_wfd_rd_7),
    .io_deq_bits_wfd_mask_0(result_v_io_deq_bits_wfd_mask_0),
    .io_deq_bits_wfd_mask_1(result_v_io_deq_bits_wfd_mask_1),
    .io_deq_bits_wfd_mask_2(result_v_io_deq_bits_wfd_mask_2),
    .io_deq_bits_wfd_mask_3(result_v_io_deq_bits_wfd_mask_3),
    .io_deq_bits_wfd_mask_4(result_v_io_deq_bits_wfd_mask_4),
    .io_deq_bits_wfd_mask_5(result_v_io_deq_bits_wfd_mask_5),
    .io_deq_bits_wfd_mask_6(result_v_io_deq_bits_wfd_mask_6),
    .io_deq_bits_wfd_mask_7(result_v_io_deq_bits_wfd_mask_7),
    .io_deq_bits_wfd(result_v_io_deq_bits_wfd),
    .io_deq_bits_reg_idxw(result_v_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_v_io_deq_bits_warp_id)
  );
  Queue_44 data_buffer ( // @[Decoupled.scala 361:21]
    .clock(data_buffer_clock),
    .reset(data_buffer_reset),
    .io_enq_ready(data_buffer_io_enq_ready),
    .io_enq_valid(data_buffer_io_enq_valid),
    .io_enq_bits_in1_0(data_buffer_io_enq_bits_in1_0),
    .io_enq_bits_in1_1(data_buffer_io_enq_bits_in1_1),
    .io_enq_bits_in1_2(data_buffer_io_enq_bits_in1_2),
    .io_enq_bits_in1_3(data_buffer_io_enq_bits_in1_3),
    .io_enq_bits_in1_4(data_buffer_io_enq_bits_in1_4),
    .io_enq_bits_in1_5(data_buffer_io_enq_bits_in1_5),
    .io_enq_bits_in1_6(data_buffer_io_enq_bits_in1_6),
    .io_enq_bits_in1_7(data_buffer_io_enq_bits_in1_7),
    .io_enq_bits_in2_0(data_buffer_io_enq_bits_in2_0),
    .io_enq_bits_in2_1(data_buffer_io_enq_bits_in2_1),
    .io_enq_bits_in2_2(data_buffer_io_enq_bits_in2_2),
    .io_enq_bits_in2_3(data_buffer_io_enq_bits_in2_3),
    .io_enq_bits_in2_4(data_buffer_io_enq_bits_in2_4),
    .io_enq_bits_in2_5(data_buffer_io_enq_bits_in2_5),
    .io_enq_bits_in2_6(data_buffer_io_enq_bits_in2_6),
    .io_enq_bits_in2_7(data_buffer_io_enq_bits_in2_7),
    .io_enq_bits_mask_0(data_buffer_io_enq_bits_mask_0),
    .io_enq_bits_mask_1(data_buffer_io_enq_bits_mask_1),
    .io_enq_bits_mask_2(data_buffer_io_enq_bits_mask_2),
    .io_enq_bits_mask_3(data_buffer_io_enq_bits_mask_3),
    .io_enq_bits_mask_4(data_buffer_io_enq_bits_mask_4),
    .io_enq_bits_mask_5(data_buffer_io_enq_bits_mask_5),
    .io_enq_bits_mask_6(data_buffer_io_enq_bits_mask_6),
    .io_enq_bits_mask_7(data_buffer_io_enq_bits_mask_7),
    .io_enq_bits_ctrl_wid(data_buffer_io_enq_bits_ctrl_wid),
    .io_enq_bits_ctrl_fp(data_buffer_io_enq_bits_ctrl_fp),
    .io_enq_bits_ctrl_reverse(data_buffer_io_enq_bits_ctrl_reverse),
    .io_enq_bits_ctrl_isvec(data_buffer_io_enq_bits_ctrl_isvec),
    .io_enq_bits_ctrl_alu_fn(data_buffer_io_enq_bits_ctrl_alu_fn),
    .io_enq_bits_ctrl_reg_idxw(data_buffer_io_enq_bits_ctrl_reg_idxw),
    .io_enq_bits_ctrl_wfd(data_buffer_io_enq_bits_ctrl_wfd),
    .io_enq_bits_ctrl_wxd(data_buffer_io_enq_bits_ctrl_wxd),
    .io_deq_ready(data_buffer_io_deq_ready),
    .io_deq_valid(data_buffer_io_deq_valid),
    .io_deq_bits_in1_0(data_buffer_io_deq_bits_in1_0),
    .io_deq_bits_in1_1(data_buffer_io_deq_bits_in1_1),
    .io_deq_bits_in1_2(data_buffer_io_deq_bits_in1_2),
    .io_deq_bits_in1_3(data_buffer_io_deq_bits_in1_3),
    .io_deq_bits_in1_4(data_buffer_io_deq_bits_in1_4),
    .io_deq_bits_in1_5(data_buffer_io_deq_bits_in1_5),
    .io_deq_bits_in1_6(data_buffer_io_deq_bits_in1_6),
    .io_deq_bits_in1_7(data_buffer_io_deq_bits_in1_7),
    .io_deq_bits_in2_0(data_buffer_io_deq_bits_in2_0),
    .io_deq_bits_in2_1(data_buffer_io_deq_bits_in2_1),
    .io_deq_bits_in2_2(data_buffer_io_deq_bits_in2_2),
    .io_deq_bits_in2_3(data_buffer_io_deq_bits_in2_3),
    .io_deq_bits_in2_4(data_buffer_io_deq_bits_in2_4),
    .io_deq_bits_in2_5(data_buffer_io_deq_bits_in2_5),
    .io_deq_bits_in2_6(data_buffer_io_deq_bits_in2_6),
    .io_deq_bits_in2_7(data_buffer_io_deq_bits_in2_7),
    .io_deq_bits_mask_0(data_buffer_io_deq_bits_mask_0),
    .io_deq_bits_mask_1(data_buffer_io_deq_bits_mask_1),
    .io_deq_bits_mask_2(data_buffer_io_deq_bits_mask_2),
    .io_deq_bits_mask_3(data_buffer_io_deq_bits_mask_3),
    .io_deq_bits_mask_4(data_buffer_io_deq_bits_mask_4),
    .io_deq_bits_mask_5(data_buffer_io_deq_bits_mask_5),
    .io_deq_bits_mask_6(data_buffer_io_deq_bits_mask_6),
    .io_deq_bits_mask_7(data_buffer_io_deq_bits_mask_7),
    .io_deq_bits_ctrl_wid(data_buffer_io_deq_bits_ctrl_wid),
    .io_deq_bits_ctrl_fp(data_buffer_io_deq_bits_ctrl_fp),
    .io_deq_bits_ctrl_reverse(data_buffer_io_deq_bits_ctrl_reverse),
    .io_deq_bits_ctrl_isvec(data_buffer_io_deq_bits_ctrl_isvec),
    .io_deq_bits_ctrl_alu_fn(data_buffer_io_deq_bits_ctrl_alu_fn),
    .io_deq_bits_ctrl_reg_idxw(data_buffer_io_deq_bits_ctrl_reg_idxw),
    .io_deq_bits_ctrl_wfd(data_buffer_io_deq_bits_ctrl_wfd),
    .io_deq_bits_ctrl_wxd(data_buffer_io_deq_bits_ctrl_wxd)
  );
  IntDivMod IntDivMod ( // @[execution.scala 209:46]
    .clock(IntDivMod_clock),
    .reset(IntDivMod_reset),
    .io_in_ready(IntDivMod_io_in_ready),
    .io_in_valid(IntDivMod_io_in_valid),
    .io_in_bits_a(IntDivMod_io_in_bits_a),
    .io_in_bits_d(IntDivMod_io_in_bits_d),
    .io_in_bits_signed(IntDivMod_io_in_bits_signed),
    .io_out_ready(IntDivMod_io_out_ready),
    .io_out_valid(IntDivMod_io_out_valid),
    .io_out_bits_q(IntDivMod_io_out_bits_q),
    .io_out_bits_r(IntDivMod_io_out_bits_r)
  );
  IntDivMod IntDivMod_1 ( // @[execution.scala 209:46]
    .clock(IntDivMod_1_clock),
    .reset(IntDivMod_1_reset),
    .io_in_ready(IntDivMod_1_io_in_ready),
    .io_in_valid(IntDivMod_1_io_in_valid),
    .io_in_bits_a(IntDivMod_1_io_in_bits_a),
    .io_in_bits_d(IntDivMod_1_io_in_bits_d),
    .io_in_bits_signed(IntDivMod_1_io_in_bits_signed),
    .io_out_ready(IntDivMod_1_io_out_ready),
    .io_out_valid(IntDivMod_1_io_out_valid),
    .io_out_bits_q(IntDivMod_1_io_out_bits_q),
    .io_out_bits_r(IntDivMod_1_io_out_bits_r)
  );
  FloatDivSqrt FloatDivSqrt ( // @[execution.scala 210:48]
    .clock(FloatDivSqrt_clock),
    .reset(FloatDivSqrt_reset),
    .io_in_ready(FloatDivSqrt_io_in_ready),
    .io_in_valid(FloatDivSqrt_io_in_valid),
    .io_in_bits_op(FloatDivSqrt_io_in_bits_op),
    .io_in_bits_a(FloatDivSqrt_io_in_bits_a),
    .io_in_bits_b(FloatDivSqrt_io_in_bits_b),
    .io_in_bits_rm(FloatDivSqrt_io_in_bits_rm),
    .io_out_ready(FloatDivSqrt_io_out_ready),
    .io_out_valid(FloatDivSqrt_io_out_valid),
    .io_out_bits_result(FloatDivSqrt_io_out_bits_result)
  );
  FloatDivSqrt FloatDivSqrt_1 ( // @[execution.scala 210:48]
    .clock(FloatDivSqrt_1_clock),
    .reset(FloatDivSqrt_1_reset),
    .io_in_ready(FloatDivSqrt_1_io_in_ready),
    .io_in_valid(FloatDivSqrt_1_io_in_valid),
    .io_in_bits_op(FloatDivSqrt_1_io_in_bits_op),
    .io_in_bits_a(FloatDivSqrt_1_io_in_bits_a),
    .io_in_bits_b(FloatDivSqrt_1_io_in_bits_b),
    .io_in_bits_rm(FloatDivSqrt_1_io_in_bits_rm),
    .io_out_ready(FloatDivSqrt_1_io_out_ready),
    .io_out_valid(FloatDivSqrt_1_io_out_valid),
    .io_out_bits_result(FloatDivSqrt_1_io_out_bits_result)
  );
  Arbiter_9 Arbiter ( // @[execution.scala 211:55]
    .io_in_0_ready(Arbiter_io_in_0_ready),
    .io_in_0_valid(Arbiter_io_in_0_valid),
    .io_in_0_bits(Arbiter_io_in_0_bits),
    .io_in_1_ready(Arbiter_io_in_1_ready),
    .io_in_1_valid(Arbiter_io_in_1_valid),
    .io_in_1_bits(Arbiter_io_in_1_bits),
    .io_out_ready(Arbiter_io_out_ready),
    .io_out_valid(Arbiter_io_out_valid),
    .io_out_bits(Arbiter_io_out_bits)
  );
  Arbiter_9 Arbiter_1 ( // @[execution.scala 211:55]
    .io_in_0_ready(Arbiter_1_io_in_0_ready),
    .io_in_0_valid(Arbiter_1_io_in_0_valid),
    .io_in_0_bits(Arbiter_1_io_in_0_bits),
    .io_in_1_ready(Arbiter_1_io_in_1_ready),
    .io_in_1_valid(Arbiter_1_io_in_1_valid),
    .io_in_1_bits(Arbiter_1_io_in_1_bits),
    .io_out_ready(Arbiter_1_io_out_ready),
    .io_out_valid(Arbiter_1_io_out_valid),
    .io_out_bits(Arbiter_1_io_out_bits)
  );
  assign io_in_ready = data_buffer_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_out_x_valid = result_x_io_deq_valid; // @[execution.scala 303:11]
  assign io_out_x_bits_wb_wxd_rd = result_x_io_deq_bits_wb_wxd_rd; // @[execution.scala 303:11]
  assign io_out_x_bits_wxd = result_x_io_deq_bits_wxd; // @[execution.scala 303:11]
  assign io_out_x_bits_reg_idxw = result_x_io_deq_bits_reg_idxw; // @[execution.scala 303:11]
  assign io_out_x_bits_warp_id = result_x_io_deq_bits_warp_id; // @[execution.scala 303:11]
  assign io_out_v_valid = result_v_io_deq_valid; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_0 = result_v_io_deq_bits_wb_wfd_rd_0; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_1 = result_v_io_deq_bits_wb_wfd_rd_1; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_2 = result_v_io_deq_bits_wb_wfd_rd_2; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_3 = result_v_io_deq_bits_wb_wfd_rd_3; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_4 = result_v_io_deq_bits_wb_wfd_rd_4; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_5 = result_v_io_deq_bits_wb_wfd_rd_5; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_6 = result_v_io_deq_bits_wb_wfd_rd_6; // @[execution.scala 302:11]
  assign io_out_v_bits_wb_wfd_rd_7 = result_v_io_deq_bits_wb_wfd_rd_7; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_0 = result_v_io_deq_bits_wfd_mask_0; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_1 = result_v_io_deq_bits_wfd_mask_1; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_2 = result_v_io_deq_bits_wfd_mask_2; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_3 = result_v_io_deq_bits_wfd_mask_3; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_4 = result_v_io_deq_bits_wfd_mask_4; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_5 = result_v_io_deq_bits_wfd_mask_5; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_6 = result_v_io_deq_bits_wfd_mask_6; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd_mask_7 = result_v_io_deq_bits_wfd_mask_7; // @[execution.scala 302:11]
  assign io_out_v_bits_wfd = result_v_io_deq_bits_wfd; // @[execution.scala 302:11]
  assign io_out_v_bits_reg_idxw = result_v_io_deq_bits_reg_idxw; // @[execution.scala 302:11]
  assign io_out_v_bits_warp_id = result_v_io_deq_bits_warp_id; // @[execution.scala 302:11]
  assign result_x_clock = clock;
  assign result_x_reset = reset;
  assign result_x_io_enq_valid = state == 2'h2 & data_buffer_io_deq_bits_ctrl_wxd; // @[execution.scala 225:42]
  assign result_x_io_enq_bits_wb_wxd_rd = out_data_0; // @[execution.scala 223:33]
  assign result_x_io_enq_bits_wxd = data_buffer_io_deq_bits_ctrl_wxd; // @[execution.scala 220:27]
  assign result_x_io_enq_bits_reg_idxw = data_buffer_io_deq_bits_ctrl_reg_idxw; // @[execution.scala 222:32]
  assign result_x_io_enq_bits_warp_id = data_buffer_io_deq_bits_ctrl_wid; // @[execution.scala 221:31]
  assign result_x_io_deq_ready = io_out_x_ready; // @[execution.scala 303:11]
  assign result_v_clock = clock;
  assign result_v_reset = reset;
  assign result_v_io_enq_valid = _result_x_io_enq_valid_T & data_buffer_io_deq_bits_ctrl_wfd; // @[execution.scala 226:42]
  assign result_v_io_enq_bits_wb_wfd_rd_0 = out_data_0; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_1 = out_data_1; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_2 = out_data_2; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_3 = out_data_3; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_4 = out_data_4; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_5 = out_data_5; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_6 = out_data_6; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wb_wfd_rd_7 = out_data_7; // @[execution.scala 217:33]
  assign result_v_io_enq_bits_wfd_mask_0 = data_buffer_io_deq_bits_mask_0; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_1 = data_buffer_io_deq_bits_mask_1; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_2 = data_buffer_io_deq_bits_mask_2; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_3 = data_buffer_io_deq_bits_mask_3; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_4 = data_buffer_io_deq_bits_mask_4; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_5 = data_buffer_io_deq_bits_mask_5; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_6 = data_buffer_io_deq_bits_mask_6; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd_mask_7 = data_buffer_io_deq_bits_mask_7; // @[execution.scala 215:32]
  assign result_v_io_enq_bits_wfd = data_buffer_io_deq_bits_ctrl_wfd; // @[execution.scala 216:27]
  assign result_v_io_enq_bits_reg_idxw = data_buffer_io_deq_bits_ctrl_reg_idxw; // @[execution.scala 218:32]
  assign result_v_io_enq_bits_warp_id = data_buffer_io_deq_bits_ctrl_wid; // @[execution.scala 219:31]
  assign result_v_io_deq_ready = io_out_v_ready; // @[execution.scala 302:11]
  assign data_buffer_clock = clock;
  assign data_buffer_reset = reset;
  assign data_buffer_io_enq_valid = io_in_valid; // @[Decoupled.scala 363:22]
  assign data_buffer_io_enq_bits_in1_0 = io_in_bits_in1_0; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_1 = io_in_bits_in1_1; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_2 = io_in_bits_in1_2; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_3 = io_in_bits_in1_3; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_4 = io_in_bits_in1_4; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_5 = io_in_bits_in1_5; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_6 = io_in_bits_in1_6; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in1_7 = io_in_bits_in1_7; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_0 = io_in_bits_in2_0; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_1 = io_in_bits_in2_1; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_2 = io_in_bits_in2_2; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_3 = io_in_bits_in2_3; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_4 = io_in_bits_in2_4; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_5 = io_in_bits_in2_5; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_6 = io_in_bits_in2_6; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_in2_7 = io_in_bits_in2_7; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_0 = io_in_bits_mask_0; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_1 = io_in_bits_mask_1; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_2 = io_in_bits_mask_2; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_3 = io_in_bits_mask_3; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_4 = io_in_bits_mask_4; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_5 = io_in_bits_mask_5; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_6 = io_in_bits_mask_6; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_mask_7 = io_in_bits_mask_7; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_wid = io_in_bits_ctrl_wid; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_fp = io_in_bits_ctrl_fp; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_reverse = io_in_bits_ctrl_reverse; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_isvec = io_in_bits_ctrl_isvec; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_alu_fn = io_in_bits_ctrl_alu_fn; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_wfd = io_in_bits_ctrl_wfd; // @[Decoupled.scala 364:21]
  assign data_buffer_io_enq_bits_ctrl_wxd = io_in_bits_ctrl_wxd; // @[Decoupled.scala 364:21]
  assign data_buffer_io_deq_ready = _result_x_io_enq_valid_T & o_ready; // @[execution.scala 257:38]
  assign IntDivMod_clock = clock;
  assign IntDivMod_reset = reset;
  assign IntDivMod_io_in_valid = ~data_buffer_io_deq_bits_ctrl_fp & i_valid; // @[execution.scala 253:38]
  assign IntDivMod_io_in_bits_a = _T_18 & i_mask_0 ? i_data1_0 : _GEN_42; // @[execution.scala 243:41 244:25]
  assign IntDivMod_io_in_bits_d = _T_18 & i_mask_0 ? i_data2_0 : _GEN_43; // @[execution.scala 243:41 245:25]
  assign IntDivMod_io_in_bits_signed = ~data_buffer_io_deq_bits_ctrl_alu_fn[1]; // @[execution.scala 249:33]
  assign IntDivMod_io_out_ready = Arbiter_io_in_0_ready; // @[execution.scala 211:{30,30}]
  assign IntDivMod_1_clock = clock;
  assign IntDivMod_1_reset = reset;
  assign IntDivMod_1_io_in_valid = ~data_buffer_io_deq_bits_ctrl_fp & i_valid; // @[execution.scala 253:38]
  assign IntDivMod_1_io_in_bits_a = _T_18 & i_mask_1 ? i_data1_1 : _GEN_62; // @[execution.scala 243:41 244:25]
  assign IntDivMod_1_io_in_bits_d = _T_18 & i_mask_1 ? i_data2_1 : _GEN_63; // @[execution.scala 243:41 245:25]
  assign IntDivMod_1_io_in_bits_signed = ~data_buffer_io_deq_bits_ctrl_alu_fn[1]; // @[execution.scala 249:33]
  assign IntDivMod_1_io_out_ready = Arbiter_1_io_in_0_ready; // @[execution.scala 211:{30,30}]
  assign FloatDivSqrt_clock = clock;
  assign FloatDivSqrt_reset = reset;
  assign FloatDivSqrt_io_in_valid = data_buffer_io_deq_bits_ctrl_fp & i_valid; // @[execution.scala 254:39]
  assign FloatDivSqrt_io_in_bits_op = data_buffer_io_deq_bits_ctrl_alu_fn[2:0]; // @[execution.scala 251:44]
  assign FloatDivSqrt_io_in_bits_a = _T_18 & i_mask_0 ? i_data1_0 : _GEN_44; // @[execution.scala 243:41 246:27]
  assign FloatDivSqrt_io_in_bits_b = _T_18 & i_mask_0 ? i_data2_0 : _GEN_45; // @[execution.scala 243:41 247:27]
  assign FloatDivSqrt_io_in_bits_rm = io_rm; // @[execution.scala 210:23 250:28]
  assign FloatDivSqrt_io_out_ready = Arbiter_io_in_1_ready; // @[execution.scala 211:{30,30}]
  assign FloatDivSqrt_1_clock = clock;
  assign FloatDivSqrt_1_reset = reset;
  assign FloatDivSqrt_1_io_in_valid = data_buffer_io_deq_bits_ctrl_fp & i_valid; // @[execution.scala 254:39]
  assign FloatDivSqrt_1_io_in_bits_op = data_buffer_io_deq_bits_ctrl_alu_fn[2:0]; // @[execution.scala 251:44]
  assign FloatDivSqrt_1_io_in_bits_a = _T_18 & i_mask_1 ? i_data1_1 : _GEN_64; // @[execution.scala 243:41 246:27]
  assign FloatDivSqrt_1_io_in_bits_b = _T_18 & i_mask_1 ? i_data2_1 : _GEN_65; // @[execution.scala 243:41 247:27]
  assign FloatDivSqrt_1_io_in_bits_rm = io_rm; // @[execution.scala 210:23 250:28]
  assign FloatDivSqrt_1_io_out_ready = Arbiter_1_io_in_1_ready; // @[execution.scala 211:{30,30}]
  assign Arbiter_io_in_0_valid = IntDivMod_io_out_valid; // @[execution.scala 209:{21,21}]
  assign Arbiter_io_in_0_bits = data_buffer_io_deq_bits_ctrl_alu_fn[0] ? intDiv_0_out_bits_r : intDiv_0_out_bits_q; // @[execution.scala 230:41]
  assign Arbiter_io_in_1_valid = FloatDivSqrt_io_out_valid; // @[execution.scala 210:{23,23}]
  assign Arbiter_io_in_1_bits = FloatDivSqrt_io_out_bits_result; // @[execution.scala 210:{23,23}]
  assign Arbiter_io_out_ready = alu_out_arbiter_0_out_valid & alu_out_arbiter_1_out_valid; // @[execution.scala 212:87]
  assign Arbiter_1_io_in_0_valid = IntDivMod_1_io_out_valid; // @[execution.scala 209:{21,21}]
  assign Arbiter_1_io_in_0_bits = data_buffer_io_deq_bits_ctrl_alu_fn[0] ? intDiv_1_out_bits_r : intDiv_1_out_bits_q; // @[execution.scala 230:41]
  assign Arbiter_1_io_in_1_valid = FloatDivSqrt_1_io_out_valid; // @[execution.scala 210:{23,23}]
  assign Arbiter_1_io_in_1_bits = FloatDivSqrt_1_io_out_bits_result; // @[execution.scala 210:{23,23}]
  assign Arbiter_1_io_out_ready = alu_out_arbiter_0_out_valid & alu_out_arbiter_1_out_valid; // @[execution.scala 212:87]
  always @(posedge clock) begin
    if (reset) begin // @[execution.scala 179:20]
      state <= 2'h0; // @[execution.scala 179:20]
    end else if (2'h0 == state) begin // @[execution.scala 260:16]
      if (_T_41) begin // @[execution.scala 262:25]
        state <= 2'h1; // @[execution.scala 263:14]
      end
    end else if (2'h1 == state) begin // @[execution.scala 260:16]
      if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
        state <= _GEN_103;
      end else begin
        state <= _GEN_105;
      end
    end else if (2'h2 == state) begin // @[execution.scala 260:16]
      state <= _GEN_118;
    end
    mask <= _GEN_163[7:0]; // @[execution.scala 182:{19,19}]
    if (reset) begin // @[execution.scala 189:23]
      out_data_0 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_0 <= _GEN_80;
        end else begin
          out_data_0 <= _GEN_104;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_0 <= _GEN_119;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_1 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_1 <= _GEN_81;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_1 <= _GEN_120;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_2 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_2 <= _GEN_87;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_2 <= _GEN_121;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_3 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_3 <= _GEN_88;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_3 <= _GEN_122;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_4 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_4 <= _GEN_94;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_4 <= _GEN_123;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_5 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_5 <= _GEN_95;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_5 <= _GEN_124;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_6 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_6 <= _GEN_101;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_6 <= _GEN_125;
      end
    end
    if (reset) begin // @[execution.scala 189:23]
      out_data_7 <= 32'h0; // @[execution.scala 189:23]
    end else if (!(2'h0 == state)) begin // @[execution.scala 260:16]
      if (2'h1 == state) begin // @[execution.scala 260:16]
        if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
          out_data_7 <= _GEN_102;
        end
      end else if (2'h2 == state) begin // @[execution.scala 260:16]
        out_data_7 <= _GEN_126;
      end
    end
    if (reset) begin // @[execution.scala 193:24]
      i_valid <= 1'h0; // @[execution.scala 193:24]
    end else if (2'h0 == state) begin // @[execution.scala 260:16]
      i_valid <= _GEN_74;
    end else if (2'h1 == state) begin // @[execution.scala 260:16]
      if (data_buffer_io_deq_bits_ctrl_isvec & alu_out_fire) begin // @[execution.scala 272:56]
        i_valid <= _GEN_100;
      end else begin
        i_valid <= _GEN_106;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  out_data_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  out_data_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  out_data_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  out_data_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  out_data_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  out_data_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  out_data_6 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  out_data_7 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  i_valid = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU2WB(
  output        io_lsu_rsp_ready,
  input         io_lsu_rsp_valid,
  input  [1:0]  io_lsu_rsp_bits_tag_warp_id,
  input         io_lsu_rsp_bits_tag_wfd,
  input         io_lsu_rsp_bits_tag_wxd,
  input  [4:0]  io_lsu_rsp_bits_tag_reg_idxw,
  input         io_lsu_rsp_bits_tag_mask_0,
  input         io_lsu_rsp_bits_tag_mask_1,
  input         io_lsu_rsp_bits_tag_mask_2,
  input         io_lsu_rsp_bits_tag_mask_3,
  input         io_lsu_rsp_bits_tag_mask_4,
  input         io_lsu_rsp_bits_tag_mask_5,
  input         io_lsu_rsp_bits_tag_mask_6,
  input         io_lsu_rsp_bits_tag_mask_7,
  input         io_lsu_rsp_bits_tag_isWrite,
  input  [31:0] io_lsu_rsp_bits_data_0,
  input  [31:0] io_lsu_rsp_bits_data_1,
  input  [31:0] io_lsu_rsp_bits_data_2,
  input  [31:0] io_lsu_rsp_bits_data_3,
  input  [31:0] io_lsu_rsp_bits_data_4,
  input  [31:0] io_lsu_rsp_bits_data_5,
  input  [31:0] io_lsu_rsp_bits_data_6,
  input  [31:0] io_lsu_rsp_bits_data_7,
  input         io_out_x_ready,
  output        io_out_x_valid,
  output [31:0] io_out_x_bits_wb_wxd_rd,
  output        io_out_x_bits_wxd,
  output [4:0]  io_out_x_bits_reg_idxw,
  output [1:0]  io_out_x_bits_warp_id,
  input         io_out_v_ready,
  output        io_out_v_valid,
  output [31:0] io_out_v_bits_wb_wfd_rd_0,
  output [31:0] io_out_v_bits_wb_wfd_rd_1,
  output [31:0] io_out_v_bits_wb_wfd_rd_2,
  output [31:0] io_out_v_bits_wb_wfd_rd_3,
  output [31:0] io_out_v_bits_wb_wfd_rd_4,
  output [31:0] io_out_v_bits_wb_wfd_rd_5,
  output [31:0] io_out_v_bits_wb_wfd_rd_6,
  output [31:0] io_out_v_bits_wb_wfd_rd_7,
  output        io_out_v_bits_wfd_mask_0,
  output        io_out_v_bits_wfd_mask_1,
  output        io_out_v_bits_wfd_mask_2,
  output        io_out_v_bits_wfd_mask_3,
  output        io_out_v_bits_wfd_mask_4,
  output        io_out_v_bits_wfd_mask_5,
  output        io_out_v_bits_wfd_mask_6,
  output        io_out_v_bits_wfd_mask_7,
  output        io_out_v_bits_wfd,
  output [4:0]  io_out_v_bits_reg_idxw,
  output [1:0]  io_out_v_bits_warp_id
);
  wire  _GEN_0 = io_lsu_rsp_bits_tag_wfd & io_lsu_rsp_valid; // @[LSU.scala 311:38 312:19 316:21]
  wire  _GEN_2 = io_lsu_rsp_bits_tag_wfd ? io_out_v_ready : io_lsu_rsp_bits_tag_isWrite; // @[LSU.scala 311:38 314:21 318:23]
  assign io_lsu_rsp_ready = io_lsu_rsp_bits_tag_wxd ? io_out_x_ready : _GEN_2; // @[LSU.scala 307:32 310:21]
  assign io_out_x_valid = io_lsu_rsp_bits_tag_wxd & io_lsu_rsp_valid; // @[LSU.scala 307:32 308:19]
  assign io_out_x_bits_wb_wxd_rd = io_lsu_rsp_bits_data_0; // @[LSU.scala 301:26]
  assign io_out_x_bits_wxd = io_lsu_rsp_bits_tag_wxd; // @[LSU.scala 300:20]
  assign io_out_x_bits_reg_idxw = io_lsu_rsp_bits_tag_reg_idxw; // @[LSU.scala 299:25]
  assign io_out_x_bits_warp_id = io_lsu_rsp_bits_tag_warp_id; // @[LSU.scala 298:24]
  assign io_out_v_valid = io_lsu_rsp_bits_tag_wxd ? 1'h0 : _GEN_0; // @[LSU.scala 307:32 309:19]
  assign io_out_v_bits_wb_wfd_rd_0 = io_lsu_rsp_bits_data_0; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_1 = io_lsu_rsp_bits_data_1; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_2 = io_lsu_rsp_bits_data_2; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_3 = io_lsu_rsp_bits_data_3; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_4 = io_lsu_rsp_bits_data_4; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_5 = io_lsu_rsp_bits_data_5; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_6 = io_lsu_rsp_bits_data_6; // @[LSU.scala 306:26]
  assign io_out_v_bits_wb_wfd_rd_7 = io_lsu_rsp_bits_data_7; // @[LSU.scala 306:26]
  assign io_out_v_bits_wfd_mask_0 = io_lsu_rsp_bits_tag_mask_0; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_1 = io_lsu_rsp_bits_tag_mask_1; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_2 = io_lsu_rsp_bits_tag_mask_2; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_3 = io_lsu_rsp_bits_tag_mask_3; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_4 = io_lsu_rsp_bits_tag_mask_4; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_5 = io_lsu_rsp_bits_tag_mask_5; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_6 = io_lsu_rsp_bits_tag_mask_6; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd_mask_7 = io_lsu_rsp_bits_tag_mask_7; // @[LSU.scala 305:25]
  assign io_out_v_bits_wfd = io_lsu_rsp_bits_tag_wfd; // @[LSU.scala 304:20]
  assign io_out_v_bits_reg_idxw = io_lsu_rsp_bits_tag_reg_idxw; // @[LSU.scala 303:25]
  assign io_out_v_bits_warp_id = io_lsu_rsp_bits_tag_warp_id; // @[LSU.scala 302:24]
endmodule
module Arbiter_11(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_wb_wxd_rd,
  input         io_in_0_bits_wxd,
  input  [4:0]  io_in_0_bits_reg_idxw,
  input  [1:0]  io_in_0_bits_warp_id,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_wb_wxd_rd,
  input         io_in_1_bits_wxd,
  input  [4:0]  io_in_1_bits_reg_idxw,
  input  [1:0]  io_in_1_bits_warp_id,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_wb_wxd_rd,
  input         io_in_2_bits_wxd,
  input  [4:0]  io_in_2_bits_reg_idxw,
  input  [1:0]  io_in_2_bits_warp_id,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_wb_wxd_rd,
  input         io_in_3_bits_wxd,
  input  [4:0]  io_in_3_bits_reg_idxw,
  input  [1:0]  io_in_3_bits_warp_id,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [31:0] io_in_4_bits_wb_wxd_rd,
  input         io_in_4_bits_wxd,
  input  [4:0]  io_in_4_bits_reg_idxw,
  input  [1:0]  io_in_4_bits_warp_id,
  output        io_out_valid,
  output [31:0] io_out_bits_wb_wxd_rd,
  output        io_out_bits_wxd,
  output [4:0]  io_out_bits_reg_idxw,
  output [1:0]  io_out_bits_warp_id
);
  wire [1:0] _GEN_1 = io_in_3_valid ? io_in_3_bits_warp_id : io_in_4_bits_warp_id; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [4:0] _GEN_2 = io_in_3_valid ? io_in_3_bits_reg_idxw : io_in_4_bits_reg_idxw; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_3 = io_in_3_valid ? io_in_3_bits_wxd : io_in_4_bits_wxd; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_4 = io_in_3_valid ? io_in_3_bits_wb_wxd_rd : io_in_4_bits_wb_wxd_rd; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [1:0] _GEN_6 = io_in_2_valid ? io_in_2_bits_warp_id : _GEN_1; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_7 = io_in_2_valid ? io_in_2_bits_reg_idxw : _GEN_2; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_8 = io_in_2_valid ? io_in_2_bits_wxd : _GEN_3; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_9 = io_in_2_valid ? io_in_2_bits_wb_wxd_rd : _GEN_4; // @[Arbiter.scala 141:26 143:19]
  wire [1:0] _GEN_11 = io_in_1_valid ? io_in_1_bits_warp_id : _GEN_6; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_12 = io_in_1_valid ? io_in_1_bits_reg_idxw : _GEN_7; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_13 = io_in_1_valid ? io_in_1_bits_wxd : _GEN_8; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_14 = io_in_1_valid ? io_in_1_bits_wb_wxd_rd : _GEN_9; // @[Arbiter.scala 141:26 143:19]
  wire  grant_4 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid); // @[Arbiter.scala 46:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 46:78]
  assign io_in_3_ready = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 46:78]
  assign io_in_4_ready = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid); // @[Arbiter.scala 46:78]
  assign io_out_valid = ~grant_4 | io_in_4_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_wb_wxd_rd = io_in_0_valid ? io_in_0_bits_wb_wxd_rd : _GEN_14; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wxd = io_in_0_valid ? io_in_0_bits_wxd : _GEN_13; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_reg_idxw = io_in_0_valid ? io_in_0_bits_reg_idxw : _GEN_12; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_warp_id = io_in_0_valid ? io_in_0_bits_warp_id : _GEN_11; // @[Arbiter.scala 141:26 143:19]
endmodule
module Arbiter_12(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_wb_wfd_rd_0,
  input  [31:0] io_in_0_bits_wb_wfd_rd_1,
  input  [31:0] io_in_0_bits_wb_wfd_rd_2,
  input  [31:0] io_in_0_bits_wb_wfd_rd_3,
  input  [31:0] io_in_0_bits_wb_wfd_rd_4,
  input  [31:0] io_in_0_bits_wb_wfd_rd_5,
  input  [31:0] io_in_0_bits_wb_wfd_rd_6,
  input  [31:0] io_in_0_bits_wb_wfd_rd_7,
  input         io_in_0_bits_wfd_mask_0,
  input         io_in_0_bits_wfd_mask_1,
  input         io_in_0_bits_wfd_mask_2,
  input         io_in_0_bits_wfd_mask_3,
  input         io_in_0_bits_wfd_mask_4,
  input         io_in_0_bits_wfd_mask_5,
  input         io_in_0_bits_wfd_mask_6,
  input         io_in_0_bits_wfd_mask_7,
  input         io_in_0_bits_wfd,
  input  [4:0]  io_in_0_bits_reg_idxw,
  input  [1:0]  io_in_0_bits_warp_id,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_wb_wfd_rd_0,
  input  [31:0] io_in_1_bits_wb_wfd_rd_1,
  input  [31:0] io_in_1_bits_wb_wfd_rd_2,
  input  [31:0] io_in_1_bits_wb_wfd_rd_3,
  input  [31:0] io_in_1_bits_wb_wfd_rd_4,
  input  [31:0] io_in_1_bits_wb_wfd_rd_5,
  input  [31:0] io_in_1_bits_wb_wfd_rd_6,
  input  [31:0] io_in_1_bits_wb_wfd_rd_7,
  input         io_in_1_bits_wfd_mask_0,
  input         io_in_1_bits_wfd_mask_1,
  input         io_in_1_bits_wfd_mask_2,
  input         io_in_1_bits_wfd_mask_3,
  input         io_in_1_bits_wfd_mask_4,
  input         io_in_1_bits_wfd_mask_5,
  input         io_in_1_bits_wfd_mask_6,
  input         io_in_1_bits_wfd_mask_7,
  input         io_in_1_bits_wfd,
  input  [4:0]  io_in_1_bits_reg_idxw,
  input  [1:0]  io_in_1_bits_warp_id,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_wb_wfd_rd_0,
  input  [31:0] io_in_2_bits_wb_wfd_rd_1,
  input  [31:0] io_in_2_bits_wb_wfd_rd_2,
  input  [31:0] io_in_2_bits_wb_wfd_rd_3,
  input  [31:0] io_in_2_bits_wb_wfd_rd_4,
  input  [31:0] io_in_2_bits_wb_wfd_rd_5,
  input  [31:0] io_in_2_bits_wb_wfd_rd_6,
  input  [31:0] io_in_2_bits_wb_wfd_rd_7,
  input         io_in_2_bits_wfd_mask_0,
  input         io_in_2_bits_wfd_mask_1,
  input         io_in_2_bits_wfd_mask_2,
  input         io_in_2_bits_wfd_mask_3,
  input         io_in_2_bits_wfd_mask_4,
  input         io_in_2_bits_wfd_mask_5,
  input         io_in_2_bits_wfd_mask_6,
  input         io_in_2_bits_wfd_mask_7,
  input         io_in_2_bits_wfd,
  input  [4:0]  io_in_2_bits_reg_idxw,
  input  [1:0]  io_in_2_bits_warp_id,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_wb_wfd_rd_0,
  input  [31:0] io_in_3_bits_wb_wfd_rd_1,
  input  [31:0] io_in_3_bits_wb_wfd_rd_2,
  input  [31:0] io_in_3_bits_wb_wfd_rd_3,
  input  [31:0] io_in_3_bits_wb_wfd_rd_4,
  input  [31:0] io_in_3_bits_wb_wfd_rd_5,
  input  [31:0] io_in_3_bits_wb_wfd_rd_6,
  input  [31:0] io_in_3_bits_wb_wfd_rd_7,
  input         io_in_3_bits_wfd_mask_0,
  input         io_in_3_bits_wfd_mask_1,
  input         io_in_3_bits_wfd_mask_2,
  input         io_in_3_bits_wfd_mask_3,
  input         io_in_3_bits_wfd_mask_4,
  input         io_in_3_bits_wfd_mask_5,
  input         io_in_3_bits_wfd_mask_6,
  input         io_in_3_bits_wfd_mask_7,
  input         io_in_3_bits_wfd,
  input  [4:0]  io_in_3_bits_reg_idxw,
  input  [1:0]  io_in_3_bits_warp_id,
  output        io_out_valid,
  output [31:0] io_out_bits_wb_wfd_rd_0,
  output [31:0] io_out_bits_wb_wfd_rd_1,
  output [31:0] io_out_bits_wb_wfd_rd_2,
  output [31:0] io_out_bits_wb_wfd_rd_3,
  output [31:0] io_out_bits_wb_wfd_rd_4,
  output [31:0] io_out_bits_wb_wfd_rd_5,
  output [31:0] io_out_bits_wb_wfd_rd_6,
  output [31:0] io_out_bits_wb_wfd_rd_7,
  output        io_out_bits_wfd_mask_0,
  output        io_out_bits_wfd_mask_1,
  output        io_out_bits_wfd_mask_2,
  output        io_out_bits_wfd_mask_3,
  output        io_out_bits_wfd_mask_4,
  output        io_out_bits_wfd_mask_5,
  output        io_out_bits_wfd_mask_6,
  output        io_out_bits_wfd_mask_7,
  output        io_out_bits_wfd,
  output [4:0]  io_out_bits_reg_idxw,
  output [1:0]  io_out_bits_warp_id
);
  wire [1:0] _GEN_1 = io_in_2_valid ? io_in_2_bits_warp_id : io_in_3_bits_warp_id; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [4:0] _GEN_2 = io_in_2_valid ? io_in_2_bits_reg_idxw : io_in_3_bits_reg_idxw; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_3 = io_in_2_valid ? io_in_2_bits_wfd : io_in_3_bits_wfd; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_4 = io_in_2_valid ? io_in_2_bits_wfd_mask_0 : io_in_3_bits_wfd_mask_0; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_5 = io_in_2_valid ? io_in_2_bits_wfd_mask_1 : io_in_3_bits_wfd_mask_1; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_6 = io_in_2_valid ? io_in_2_bits_wfd_mask_2 : io_in_3_bits_wfd_mask_2; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_7 = io_in_2_valid ? io_in_2_bits_wfd_mask_3 : io_in_3_bits_wfd_mask_3; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_8 = io_in_2_valid ? io_in_2_bits_wfd_mask_4 : io_in_3_bits_wfd_mask_4; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_9 = io_in_2_valid ? io_in_2_bits_wfd_mask_5 : io_in_3_bits_wfd_mask_5; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_10 = io_in_2_valid ? io_in_2_bits_wfd_mask_6 : io_in_3_bits_wfd_mask_6; // @[Arbiter.scala 139:15 141:26 143:19]
  wire  _GEN_11 = io_in_2_valid ? io_in_2_bits_wfd_mask_7 : io_in_3_bits_wfd_mask_7; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_12 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_0 : io_in_3_bits_wb_wfd_rd_0; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_13 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_1 : io_in_3_bits_wb_wfd_rd_1; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_14 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_2 : io_in_3_bits_wb_wfd_rd_2; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_15 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_3 : io_in_3_bits_wb_wfd_rd_3; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_16 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_4 : io_in_3_bits_wb_wfd_rd_4; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_17 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_5 : io_in_3_bits_wb_wfd_rd_5; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_18 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_6 : io_in_3_bits_wb_wfd_rd_6; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_19 = io_in_2_valid ? io_in_2_bits_wb_wfd_rd_7 : io_in_3_bits_wb_wfd_rd_7; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [1:0] _GEN_21 = io_in_1_valid ? io_in_1_bits_warp_id : _GEN_1; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_22 = io_in_1_valid ? io_in_1_bits_reg_idxw : _GEN_2; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_23 = io_in_1_valid ? io_in_1_bits_wfd : _GEN_3; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_24 = io_in_1_valid ? io_in_1_bits_wfd_mask_0 : _GEN_4; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_25 = io_in_1_valid ? io_in_1_bits_wfd_mask_1 : _GEN_5; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_26 = io_in_1_valid ? io_in_1_bits_wfd_mask_2 : _GEN_6; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_27 = io_in_1_valid ? io_in_1_bits_wfd_mask_3 : _GEN_7; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_28 = io_in_1_valid ? io_in_1_bits_wfd_mask_4 : _GEN_8; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_29 = io_in_1_valid ? io_in_1_bits_wfd_mask_5 : _GEN_9; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_30 = io_in_1_valid ? io_in_1_bits_wfd_mask_6 : _GEN_10; // @[Arbiter.scala 141:26 143:19]
  wire  _GEN_31 = io_in_1_valid ? io_in_1_bits_wfd_mask_7 : _GEN_11; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_32 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_0 : _GEN_12; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_33 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_1 : _GEN_13; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_34 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_2 : _GEN_14; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_35 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_3 : _GEN_15; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_36 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_4 : _GEN_16; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_37 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_5 : _GEN_17; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_38 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_6 : _GEN_18; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_39 = io_in_1_valid ? io_in_1_bits_wb_wfd_rd_7 : _GEN_19; // @[Arbiter.scala 141:26 143:19]
  wire  grant_3 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 46:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 46:78]
  assign io_in_3_ready = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 46:78]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_wb_wfd_rd_0 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_0 : _GEN_32; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_1 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_1 : _GEN_33; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_2 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_2 : _GEN_34; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_3 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_3 : _GEN_35; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_4 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_4 : _GEN_36; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_5 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_5 : _GEN_37; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_6 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_6 : _GEN_38; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wb_wfd_rd_7 = io_in_0_valid ? io_in_0_bits_wb_wfd_rd_7 : _GEN_39; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_0 = io_in_0_valid ? io_in_0_bits_wfd_mask_0 : _GEN_24; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_1 = io_in_0_valid ? io_in_0_bits_wfd_mask_1 : _GEN_25; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_2 = io_in_0_valid ? io_in_0_bits_wfd_mask_2 : _GEN_26; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_3 = io_in_0_valid ? io_in_0_bits_wfd_mask_3 : _GEN_27; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_4 = io_in_0_valid ? io_in_0_bits_wfd_mask_4 : _GEN_28; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_5 = io_in_0_valid ? io_in_0_bits_wfd_mask_5 : _GEN_29; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_6 = io_in_0_valid ? io_in_0_bits_wfd_mask_6 : _GEN_30; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd_mask_7 = io_in_0_valid ? io_in_0_bits_wfd_mask_7 : _GEN_31; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_wfd = io_in_0_valid ? io_in_0_bits_wfd : _GEN_23; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_reg_idxw = io_in_0_valid ? io_in_0_bits_reg_idxw : _GEN_22; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_warp_id = io_in_0_valid ? io_in_0_bits_warp_id : _GEN_21; // @[Arbiter.scala 141:26 143:19]
endmodule
module Writeback(
  input         io_out_v_ready,
  output        io_out_v_valid,
  output [31:0] io_out_v_bits_wb_wfd_rd_0,
  output [31:0] io_out_v_bits_wb_wfd_rd_1,
  output [31:0] io_out_v_bits_wb_wfd_rd_2,
  output [31:0] io_out_v_bits_wb_wfd_rd_3,
  output [31:0] io_out_v_bits_wb_wfd_rd_4,
  output [31:0] io_out_v_bits_wb_wfd_rd_5,
  output [31:0] io_out_v_bits_wb_wfd_rd_6,
  output [31:0] io_out_v_bits_wb_wfd_rd_7,
  output        io_out_v_bits_wfd_mask_0,
  output        io_out_v_bits_wfd_mask_1,
  output        io_out_v_bits_wfd_mask_2,
  output        io_out_v_bits_wfd_mask_3,
  output        io_out_v_bits_wfd_mask_4,
  output        io_out_v_bits_wfd_mask_5,
  output        io_out_v_bits_wfd_mask_6,
  output        io_out_v_bits_wfd_mask_7,
  output        io_out_v_bits_wfd,
  output [4:0]  io_out_v_bits_reg_idxw,
  output [1:0]  io_out_v_bits_warp_id,
  input         io_out_x_ready,
  output        io_out_x_valid,
  output [31:0] io_out_x_bits_wb_wxd_rd,
  output        io_out_x_bits_wxd,
  output [4:0]  io_out_x_bits_reg_idxw,
  output [1:0]  io_out_x_bits_warp_id,
  input         io_in_x_0_valid,
  input  [31:0] io_in_x_0_bits_wb_wxd_rd,
  input         io_in_x_0_bits_wxd,
  input  [4:0]  io_in_x_0_bits_reg_idxw,
  input  [1:0]  io_in_x_0_bits_warp_id,
  output        io_in_x_1_ready,
  input         io_in_x_1_valid,
  input  [31:0] io_in_x_1_bits_wb_wxd_rd,
  input         io_in_x_1_bits_wxd,
  input  [4:0]  io_in_x_1_bits_reg_idxw,
  input  [1:0]  io_in_x_1_bits_warp_id,
  output        io_in_x_2_ready,
  input         io_in_x_2_valid,
  input  [31:0] io_in_x_2_bits_wb_wxd_rd,
  input         io_in_x_2_bits_wxd,
  input  [4:0]  io_in_x_2_bits_reg_idxw,
  input  [1:0]  io_in_x_2_bits_warp_id,
  output        io_in_x_3_ready,
  input         io_in_x_3_valid,
  input  [31:0] io_in_x_3_bits_wb_wxd_rd,
  input         io_in_x_3_bits_wxd,
  input  [4:0]  io_in_x_3_bits_reg_idxw,
  input  [1:0]  io_in_x_3_bits_warp_id,
  output        io_in_x_4_ready,
  input         io_in_x_4_valid,
  input  [31:0] io_in_x_4_bits_wb_wxd_rd,
  input         io_in_x_4_bits_wxd,
  input  [4:0]  io_in_x_4_bits_reg_idxw,
  input  [1:0]  io_in_x_4_bits_warp_id,
  input         io_in_v_0_valid,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_0,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_1,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_2,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_3,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_4,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_5,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_6,
  input  [31:0] io_in_v_0_bits_wb_wfd_rd_7,
  input         io_in_v_0_bits_wfd_mask_0,
  input         io_in_v_0_bits_wfd_mask_1,
  input         io_in_v_0_bits_wfd_mask_2,
  input         io_in_v_0_bits_wfd_mask_3,
  input         io_in_v_0_bits_wfd_mask_4,
  input         io_in_v_0_bits_wfd_mask_5,
  input         io_in_v_0_bits_wfd_mask_6,
  input         io_in_v_0_bits_wfd_mask_7,
  input         io_in_v_0_bits_wfd,
  input  [4:0]  io_in_v_0_bits_reg_idxw,
  input  [1:0]  io_in_v_0_bits_warp_id,
  output        io_in_v_1_ready,
  input         io_in_v_1_valid,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_0,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_1,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_2,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_3,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_4,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_5,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_6,
  input  [31:0] io_in_v_1_bits_wb_wfd_rd_7,
  input         io_in_v_1_bits_wfd_mask_0,
  input         io_in_v_1_bits_wfd_mask_1,
  input         io_in_v_1_bits_wfd_mask_2,
  input         io_in_v_1_bits_wfd_mask_3,
  input         io_in_v_1_bits_wfd_mask_4,
  input         io_in_v_1_bits_wfd_mask_5,
  input         io_in_v_1_bits_wfd_mask_6,
  input         io_in_v_1_bits_wfd_mask_7,
  input         io_in_v_1_bits_wfd,
  input  [4:0]  io_in_v_1_bits_reg_idxw,
  input  [1:0]  io_in_v_1_bits_warp_id,
  output        io_in_v_2_ready,
  input         io_in_v_2_valid,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_0,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_1,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_2,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_3,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_4,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_5,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_6,
  input  [31:0] io_in_v_2_bits_wb_wfd_rd_7,
  input         io_in_v_2_bits_wfd_mask_0,
  input         io_in_v_2_bits_wfd_mask_1,
  input         io_in_v_2_bits_wfd_mask_2,
  input         io_in_v_2_bits_wfd_mask_3,
  input         io_in_v_2_bits_wfd_mask_4,
  input         io_in_v_2_bits_wfd_mask_5,
  input         io_in_v_2_bits_wfd_mask_6,
  input         io_in_v_2_bits_wfd_mask_7,
  input         io_in_v_2_bits_wfd,
  input  [4:0]  io_in_v_2_bits_reg_idxw,
  input  [1:0]  io_in_v_2_bits_warp_id,
  output        io_in_v_3_ready,
  input         io_in_v_3_valid,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_0,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_1,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_2,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_3,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_4,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_5,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_6,
  input  [31:0] io_in_v_3_bits_wb_wfd_rd_7,
  input         io_in_v_3_bits_wfd_mask_0,
  input         io_in_v_3_bits_wfd_mask_1,
  input         io_in_v_3_bits_wfd_mask_2,
  input         io_in_v_3_bits_wfd_mask_3,
  input         io_in_v_3_bits_wfd_mask_4,
  input         io_in_v_3_bits_wfd_mask_5,
  input         io_in_v_3_bits_wfd_mask_6,
  input         io_in_v_3_bits_wfd_mask_7,
  input         io_in_v_3_bits_wfd,
  input  [4:0]  io_in_v_3_bits_reg_idxw,
  input  [1:0]  io_in_v_3_bits_warp_id
);
  wire  arbiter_x_io_in_0_valid; // @[writeback.scala 35:23]
  wire [31:0] arbiter_x_io_in_0_bits_wb_wxd_rd; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_0_bits_wxd; // @[writeback.scala 35:23]
  wire [4:0] arbiter_x_io_in_0_bits_reg_idxw; // @[writeback.scala 35:23]
  wire [1:0] arbiter_x_io_in_0_bits_warp_id; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_1_ready; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_1_valid; // @[writeback.scala 35:23]
  wire [31:0] arbiter_x_io_in_1_bits_wb_wxd_rd; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_1_bits_wxd; // @[writeback.scala 35:23]
  wire [4:0] arbiter_x_io_in_1_bits_reg_idxw; // @[writeback.scala 35:23]
  wire [1:0] arbiter_x_io_in_1_bits_warp_id; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_2_ready; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_2_valid; // @[writeback.scala 35:23]
  wire [31:0] arbiter_x_io_in_2_bits_wb_wxd_rd; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_2_bits_wxd; // @[writeback.scala 35:23]
  wire [4:0] arbiter_x_io_in_2_bits_reg_idxw; // @[writeback.scala 35:23]
  wire [1:0] arbiter_x_io_in_2_bits_warp_id; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_3_ready; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_3_valid; // @[writeback.scala 35:23]
  wire [31:0] arbiter_x_io_in_3_bits_wb_wxd_rd; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_3_bits_wxd; // @[writeback.scala 35:23]
  wire [4:0] arbiter_x_io_in_3_bits_reg_idxw; // @[writeback.scala 35:23]
  wire [1:0] arbiter_x_io_in_3_bits_warp_id; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_4_ready; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_4_valid; // @[writeback.scala 35:23]
  wire [31:0] arbiter_x_io_in_4_bits_wb_wxd_rd; // @[writeback.scala 35:23]
  wire  arbiter_x_io_in_4_bits_wxd; // @[writeback.scala 35:23]
  wire [4:0] arbiter_x_io_in_4_bits_reg_idxw; // @[writeback.scala 35:23]
  wire [1:0] arbiter_x_io_in_4_bits_warp_id; // @[writeback.scala 35:23]
  wire  arbiter_x_io_out_valid; // @[writeback.scala 35:23]
  wire [31:0] arbiter_x_io_out_bits_wb_wxd_rd; // @[writeback.scala 35:23]
  wire  arbiter_x_io_out_bits_wxd; // @[writeback.scala 35:23]
  wire [4:0] arbiter_x_io_out_bits_reg_idxw; // @[writeback.scala 35:23]
  wire [1:0] arbiter_x_io_out_bits_warp_id; // @[writeback.scala 35:23]
  wire  arbiter_v_io_in_0_valid; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_0; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_1; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_2; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_3; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_4; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_5; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_6; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_0_bits_wb_wfd_rd_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_0; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_1; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_2; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_3; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_4; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_5; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_6; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd_mask_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_0_bits_wfd; // @[writeback.scala 36:23]
  wire [4:0] arbiter_v_io_in_0_bits_reg_idxw; // @[writeback.scala 36:23]
  wire [1:0] arbiter_v_io_in_0_bits_warp_id; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_ready; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_valid; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_0; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_1; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_2; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_3; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_4; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_5; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_6; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_1_bits_wb_wfd_rd_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_0; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_1; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_2; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_3; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_4; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_5; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_6; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd_mask_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_1_bits_wfd; // @[writeback.scala 36:23]
  wire [4:0] arbiter_v_io_in_1_bits_reg_idxw; // @[writeback.scala 36:23]
  wire [1:0] arbiter_v_io_in_1_bits_warp_id; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_ready; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_valid; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_0; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_1; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_2; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_3; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_4; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_5; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_6; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_2_bits_wb_wfd_rd_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_0; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_1; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_2; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_3; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_4; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_5; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_6; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd_mask_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_2_bits_wfd; // @[writeback.scala 36:23]
  wire [4:0] arbiter_v_io_in_2_bits_reg_idxw; // @[writeback.scala 36:23]
  wire [1:0] arbiter_v_io_in_2_bits_warp_id; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_ready; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_valid; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_0; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_1; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_2; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_3; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_4; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_5; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_6; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_in_3_bits_wb_wfd_rd_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_0; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_1; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_2; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_3; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_4; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_5; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_6; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd_mask_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_in_3_bits_wfd; // @[writeback.scala 36:23]
  wire [4:0] arbiter_v_io_in_3_bits_reg_idxw; // @[writeback.scala 36:23]
  wire [1:0] arbiter_v_io_in_3_bits_warp_id; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_valid; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_0; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_1; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_2; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_3; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_4; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_5; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_6; // @[writeback.scala 36:23]
  wire [31:0] arbiter_v_io_out_bits_wb_wfd_rd_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_0; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_1; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_2; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_3; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_4; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_5; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_6; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd_mask_7; // @[writeback.scala 36:23]
  wire  arbiter_v_io_out_bits_wfd; // @[writeback.scala 36:23]
  wire [4:0] arbiter_v_io_out_bits_reg_idxw; // @[writeback.scala 36:23]
  wire [1:0] arbiter_v_io_out_bits_warp_id; // @[writeback.scala 36:23]
  Arbiter_11 arbiter_x ( // @[writeback.scala 35:23]
    .io_in_0_valid(arbiter_x_io_in_0_valid),
    .io_in_0_bits_wb_wxd_rd(arbiter_x_io_in_0_bits_wb_wxd_rd),
    .io_in_0_bits_wxd(arbiter_x_io_in_0_bits_wxd),
    .io_in_0_bits_reg_idxw(arbiter_x_io_in_0_bits_reg_idxw),
    .io_in_0_bits_warp_id(arbiter_x_io_in_0_bits_warp_id),
    .io_in_1_ready(arbiter_x_io_in_1_ready),
    .io_in_1_valid(arbiter_x_io_in_1_valid),
    .io_in_1_bits_wb_wxd_rd(arbiter_x_io_in_1_bits_wb_wxd_rd),
    .io_in_1_bits_wxd(arbiter_x_io_in_1_bits_wxd),
    .io_in_1_bits_reg_idxw(arbiter_x_io_in_1_bits_reg_idxw),
    .io_in_1_bits_warp_id(arbiter_x_io_in_1_bits_warp_id),
    .io_in_2_ready(arbiter_x_io_in_2_ready),
    .io_in_2_valid(arbiter_x_io_in_2_valid),
    .io_in_2_bits_wb_wxd_rd(arbiter_x_io_in_2_bits_wb_wxd_rd),
    .io_in_2_bits_wxd(arbiter_x_io_in_2_bits_wxd),
    .io_in_2_bits_reg_idxw(arbiter_x_io_in_2_bits_reg_idxw),
    .io_in_2_bits_warp_id(arbiter_x_io_in_2_bits_warp_id),
    .io_in_3_ready(arbiter_x_io_in_3_ready),
    .io_in_3_valid(arbiter_x_io_in_3_valid),
    .io_in_3_bits_wb_wxd_rd(arbiter_x_io_in_3_bits_wb_wxd_rd),
    .io_in_3_bits_wxd(arbiter_x_io_in_3_bits_wxd),
    .io_in_3_bits_reg_idxw(arbiter_x_io_in_3_bits_reg_idxw),
    .io_in_3_bits_warp_id(arbiter_x_io_in_3_bits_warp_id),
    .io_in_4_ready(arbiter_x_io_in_4_ready),
    .io_in_4_valid(arbiter_x_io_in_4_valid),
    .io_in_4_bits_wb_wxd_rd(arbiter_x_io_in_4_bits_wb_wxd_rd),
    .io_in_4_bits_wxd(arbiter_x_io_in_4_bits_wxd),
    .io_in_4_bits_reg_idxw(arbiter_x_io_in_4_bits_reg_idxw),
    .io_in_4_bits_warp_id(arbiter_x_io_in_4_bits_warp_id),
    .io_out_valid(arbiter_x_io_out_valid),
    .io_out_bits_wb_wxd_rd(arbiter_x_io_out_bits_wb_wxd_rd),
    .io_out_bits_wxd(arbiter_x_io_out_bits_wxd),
    .io_out_bits_reg_idxw(arbiter_x_io_out_bits_reg_idxw),
    .io_out_bits_warp_id(arbiter_x_io_out_bits_warp_id)
  );
  Arbiter_12 arbiter_v ( // @[writeback.scala 36:23]
    .io_in_0_valid(arbiter_v_io_in_0_valid),
    .io_in_0_bits_wb_wfd_rd_0(arbiter_v_io_in_0_bits_wb_wfd_rd_0),
    .io_in_0_bits_wb_wfd_rd_1(arbiter_v_io_in_0_bits_wb_wfd_rd_1),
    .io_in_0_bits_wb_wfd_rd_2(arbiter_v_io_in_0_bits_wb_wfd_rd_2),
    .io_in_0_bits_wb_wfd_rd_3(arbiter_v_io_in_0_bits_wb_wfd_rd_3),
    .io_in_0_bits_wb_wfd_rd_4(arbiter_v_io_in_0_bits_wb_wfd_rd_4),
    .io_in_0_bits_wb_wfd_rd_5(arbiter_v_io_in_0_bits_wb_wfd_rd_5),
    .io_in_0_bits_wb_wfd_rd_6(arbiter_v_io_in_0_bits_wb_wfd_rd_6),
    .io_in_0_bits_wb_wfd_rd_7(arbiter_v_io_in_0_bits_wb_wfd_rd_7),
    .io_in_0_bits_wfd_mask_0(arbiter_v_io_in_0_bits_wfd_mask_0),
    .io_in_0_bits_wfd_mask_1(arbiter_v_io_in_0_bits_wfd_mask_1),
    .io_in_0_bits_wfd_mask_2(arbiter_v_io_in_0_bits_wfd_mask_2),
    .io_in_0_bits_wfd_mask_3(arbiter_v_io_in_0_bits_wfd_mask_3),
    .io_in_0_bits_wfd_mask_4(arbiter_v_io_in_0_bits_wfd_mask_4),
    .io_in_0_bits_wfd_mask_5(arbiter_v_io_in_0_bits_wfd_mask_5),
    .io_in_0_bits_wfd_mask_6(arbiter_v_io_in_0_bits_wfd_mask_6),
    .io_in_0_bits_wfd_mask_7(arbiter_v_io_in_0_bits_wfd_mask_7),
    .io_in_0_bits_wfd(arbiter_v_io_in_0_bits_wfd),
    .io_in_0_bits_reg_idxw(arbiter_v_io_in_0_bits_reg_idxw),
    .io_in_0_bits_warp_id(arbiter_v_io_in_0_bits_warp_id),
    .io_in_1_ready(arbiter_v_io_in_1_ready),
    .io_in_1_valid(arbiter_v_io_in_1_valid),
    .io_in_1_bits_wb_wfd_rd_0(arbiter_v_io_in_1_bits_wb_wfd_rd_0),
    .io_in_1_bits_wb_wfd_rd_1(arbiter_v_io_in_1_bits_wb_wfd_rd_1),
    .io_in_1_bits_wb_wfd_rd_2(arbiter_v_io_in_1_bits_wb_wfd_rd_2),
    .io_in_1_bits_wb_wfd_rd_3(arbiter_v_io_in_1_bits_wb_wfd_rd_3),
    .io_in_1_bits_wb_wfd_rd_4(arbiter_v_io_in_1_bits_wb_wfd_rd_4),
    .io_in_1_bits_wb_wfd_rd_5(arbiter_v_io_in_1_bits_wb_wfd_rd_5),
    .io_in_1_bits_wb_wfd_rd_6(arbiter_v_io_in_1_bits_wb_wfd_rd_6),
    .io_in_1_bits_wb_wfd_rd_7(arbiter_v_io_in_1_bits_wb_wfd_rd_7),
    .io_in_1_bits_wfd_mask_0(arbiter_v_io_in_1_bits_wfd_mask_0),
    .io_in_1_bits_wfd_mask_1(arbiter_v_io_in_1_bits_wfd_mask_1),
    .io_in_1_bits_wfd_mask_2(arbiter_v_io_in_1_bits_wfd_mask_2),
    .io_in_1_bits_wfd_mask_3(arbiter_v_io_in_1_bits_wfd_mask_3),
    .io_in_1_bits_wfd_mask_4(arbiter_v_io_in_1_bits_wfd_mask_4),
    .io_in_1_bits_wfd_mask_5(arbiter_v_io_in_1_bits_wfd_mask_5),
    .io_in_1_bits_wfd_mask_6(arbiter_v_io_in_1_bits_wfd_mask_6),
    .io_in_1_bits_wfd_mask_7(arbiter_v_io_in_1_bits_wfd_mask_7),
    .io_in_1_bits_wfd(arbiter_v_io_in_1_bits_wfd),
    .io_in_1_bits_reg_idxw(arbiter_v_io_in_1_bits_reg_idxw),
    .io_in_1_bits_warp_id(arbiter_v_io_in_1_bits_warp_id),
    .io_in_2_ready(arbiter_v_io_in_2_ready),
    .io_in_2_valid(arbiter_v_io_in_2_valid),
    .io_in_2_bits_wb_wfd_rd_0(arbiter_v_io_in_2_bits_wb_wfd_rd_0),
    .io_in_2_bits_wb_wfd_rd_1(arbiter_v_io_in_2_bits_wb_wfd_rd_1),
    .io_in_2_bits_wb_wfd_rd_2(arbiter_v_io_in_2_bits_wb_wfd_rd_2),
    .io_in_2_bits_wb_wfd_rd_3(arbiter_v_io_in_2_bits_wb_wfd_rd_3),
    .io_in_2_bits_wb_wfd_rd_4(arbiter_v_io_in_2_bits_wb_wfd_rd_4),
    .io_in_2_bits_wb_wfd_rd_5(arbiter_v_io_in_2_bits_wb_wfd_rd_5),
    .io_in_2_bits_wb_wfd_rd_6(arbiter_v_io_in_2_bits_wb_wfd_rd_6),
    .io_in_2_bits_wb_wfd_rd_7(arbiter_v_io_in_2_bits_wb_wfd_rd_7),
    .io_in_2_bits_wfd_mask_0(arbiter_v_io_in_2_bits_wfd_mask_0),
    .io_in_2_bits_wfd_mask_1(arbiter_v_io_in_2_bits_wfd_mask_1),
    .io_in_2_bits_wfd_mask_2(arbiter_v_io_in_2_bits_wfd_mask_2),
    .io_in_2_bits_wfd_mask_3(arbiter_v_io_in_2_bits_wfd_mask_3),
    .io_in_2_bits_wfd_mask_4(arbiter_v_io_in_2_bits_wfd_mask_4),
    .io_in_2_bits_wfd_mask_5(arbiter_v_io_in_2_bits_wfd_mask_5),
    .io_in_2_bits_wfd_mask_6(arbiter_v_io_in_2_bits_wfd_mask_6),
    .io_in_2_bits_wfd_mask_7(arbiter_v_io_in_2_bits_wfd_mask_7),
    .io_in_2_bits_wfd(arbiter_v_io_in_2_bits_wfd),
    .io_in_2_bits_reg_idxw(arbiter_v_io_in_2_bits_reg_idxw),
    .io_in_2_bits_warp_id(arbiter_v_io_in_2_bits_warp_id),
    .io_in_3_ready(arbiter_v_io_in_3_ready),
    .io_in_3_valid(arbiter_v_io_in_3_valid),
    .io_in_3_bits_wb_wfd_rd_0(arbiter_v_io_in_3_bits_wb_wfd_rd_0),
    .io_in_3_bits_wb_wfd_rd_1(arbiter_v_io_in_3_bits_wb_wfd_rd_1),
    .io_in_3_bits_wb_wfd_rd_2(arbiter_v_io_in_3_bits_wb_wfd_rd_2),
    .io_in_3_bits_wb_wfd_rd_3(arbiter_v_io_in_3_bits_wb_wfd_rd_3),
    .io_in_3_bits_wb_wfd_rd_4(arbiter_v_io_in_3_bits_wb_wfd_rd_4),
    .io_in_3_bits_wb_wfd_rd_5(arbiter_v_io_in_3_bits_wb_wfd_rd_5),
    .io_in_3_bits_wb_wfd_rd_6(arbiter_v_io_in_3_bits_wb_wfd_rd_6),
    .io_in_3_bits_wb_wfd_rd_7(arbiter_v_io_in_3_bits_wb_wfd_rd_7),
    .io_in_3_bits_wfd_mask_0(arbiter_v_io_in_3_bits_wfd_mask_0),
    .io_in_3_bits_wfd_mask_1(arbiter_v_io_in_3_bits_wfd_mask_1),
    .io_in_3_bits_wfd_mask_2(arbiter_v_io_in_3_bits_wfd_mask_2),
    .io_in_3_bits_wfd_mask_3(arbiter_v_io_in_3_bits_wfd_mask_3),
    .io_in_3_bits_wfd_mask_4(arbiter_v_io_in_3_bits_wfd_mask_4),
    .io_in_3_bits_wfd_mask_5(arbiter_v_io_in_3_bits_wfd_mask_5),
    .io_in_3_bits_wfd_mask_6(arbiter_v_io_in_3_bits_wfd_mask_6),
    .io_in_3_bits_wfd_mask_7(arbiter_v_io_in_3_bits_wfd_mask_7),
    .io_in_3_bits_wfd(arbiter_v_io_in_3_bits_wfd),
    .io_in_3_bits_reg_idxw(arbiter_v_io_in_3_bits_reg_idxw),
    .io_in_3_bits_warp_id(arbiter_v_io_in_3_bits_warp_id),
    .io_out_valid(arbiter_v_io_out_valid),
    .io_out_bits_wb_wfd_rd_0(arbiter_v_io_out_bits_wb_wfd_rd_0),
    .io_out_bits_wb_wfd_rd_1(arbiter_v_io_out_bits_wb_wfd_rd_1),
    .io_out_bits_wb_wfd_rd_2(arbiter_v_io_out_bits_wb_wfd_rd_2),
    .io_out_bits_wb_wfd_rd_3(arbiter_v_io_out_bits_wb_wfd_rd_3),
    .io_out_bits_wb_wfd_rd_4(arbiter_v_io_out_bits_wb_wfd_rd_4),
    .io_out_bits_wb_wfd_rd_5(arbiter_v_io_out_bits_wb_wfd_rd_5),
    .io_out_bits_wb_wfd_rd_6(arbiter_v_io_out_bits_wb_wfd_rd_6),
    .io_out_bits_wb_wfd_rd_7(arbiter_v_io_out_bits_wb_wfd_rd_7),
    .io_out_bits_wfd_mask_0(arbiter_v_io_out_bits_wfd_mask_0),
    .io_out_bits_wfd_mask_1(arbiter_v_io_out_bits_wfd_mask_1),
    .io_out_bits_wfd_mask_2(arbiter_v_io_out_bits_wfd_mask_2),
    .io_out_bits_wfd_mask_3(arbiter_v_io_out_bits_wfd_mask_3),
    .io_out_bits_wfd_mask_4(arbiter_v_io_out_bits_wfd_mask_4),
    .io_out_bits_wfd_mask_5(arbiter_v_io_out_bits_wfd_mask_5),
    .io_out_bits_wfd_mask_6(arbiter_v_io_out_bits_wfd_mask_6),
    .io_out_bits_wfd_mask_7(arbiter_v_io_out_bits_wfd_mask_7),
    .io_out_bits_wfd(arbiter_v_io_out_bits_wfd),
    .io_out_bits_reg_idxw(arbiter_v_io_out_bits_reg_idxw),
    .io_out_bits_warp_id(arbiter_v_io_out_bits_warp_id)
  );
  assign io_out_v_valid = arbiter_v_io_out_valid; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_0 = arbiter_v_io_out_bits_wb_wfd_rd_0; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_1 = arbiter_v_io_out_bits_wb_wfd_rd_1; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_2 = arbiter_v_io_out_bits_wb_wfd_rd_2; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_3 = arbiter_v_io_out_bits_wb_wfd_rd_3; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_4 = arbiter_v_io_out_bits_wb_wfd_rd_4; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_5 = arbiter_v_io_out_bits_wb_wfd_rd_5; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_6 = arbiter_v_io_out_bits_wb_wfd_rd_6; // @[writeback.scala 40:19]
  assign io_out_v_bits_wb_wfd_rd_7 = arbiter_v_io_out_bits_wb_wfd_rd_7; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_0 = arbiter_v_io_out_bits_wfd_mask_0; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_1 = arbiter_v_io_out_bits_wfd_mask_1; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_2 = arbiter_v_io_out_bits_wfd_mask_2; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_3 = arbiter_v_io_out_bits_wfd_mask_3; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_4 = arbiter_v_io_out_bits_wfd_mask_4; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_5 = arbiter_v_io_out_bits_wfd_mask_5; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_6 = arbiter_v_io_out_bits_wfd_mask_6; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd_mask_7 = arbiter_v_io_out_bits_wfd_mask_7; // @[writeback.scala 40:19]
  assign io_out_v_bits_wfd = arbiter_v_io_out_bits_wfd; // @[writeback.scala 40:19]
  assign io_out_v_bits_reg_idxw = arbiter_v_io_out_bits_reg_idxw; // @[writeback.scala 40:19]
  assign io_out_v_bits_warp_id = arbiter_v_io_out_bits_warp_id; // @[writeback.scala 40:19]
  assign io_out_x_valid = arbiter_x_io_out_valid; // @[writeback.scala 39:19]
  assign io_out_x_bits_wb_wxd_rd = arbiter_x_io_out_bits_wb_wxd_rd; // @[writeback.scala 39:19]
  assign io_out_x_bits_wxd = arbiter_x_io_out_bits_wxd; // @[writeback.scala 39:19]
  assign io_out_x_bits_reg_idxw = arbiter_x_io_out_bits_reg_idxw; // @[writeback.scala 39:19]
  assign io_out_x_bits_warp_id = arbiter_x_io_out_bits_warp_id; // @[writeback.scala 39:19]
  assign io_in_x_1_ready = arbiter_x_io_in_1_ready; // @[Decoupled.scala 355:21 writeback.scala 37:18]
  assign io_in_x_2_ready = arbiter_x_io_in_2_ready; // @[Decoupled.scala 355:21 writeback.scala 37:18]
  assign io_in_x_3_ready = arbiter_x_io_in_3_ready; // @[Decoupled.scala 355:21 writeback.scala 37:18]
  assign io_in_x_4_ready = arbiter_x_io_in_4_ready; // @[Decoupled.scala 355:21 writeback.scala 37:18]
  assign io_in_v_1_ready = arbiter_v_io_in_1_ready; // @[Decoupled.scala 355:21 writeback.scala 38:18]
  assign io_in_v_2_ready = arbiter_v_io_in_2_ready; // @[Decoupled.scala 355:21 writeback.scala 38:18]
  assign io_in_v_3_ready = arbiter_v_io_in_3_ready; // @[Decoupled.scala 355:21 writeback.scala 38:18]
  assign arbiter_x_io_in_0_valid = io_in_x_0_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_x_io_in_0_bits_wb_wxd_rd = io_in_x_0_bits_wb_wxd_rd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_0_bits_wxd = io_in_x_0_bits_wxd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_0_bits_reg_idxw = io_in_x_0_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_0_bits_warp_id = io_in_x_0_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_1_valid = io_in_x_1_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_x_io_in_1_bits_wb_wxd_rd = io_in_x_1_bits_wb_wxd_rd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_1_bits_wxd = io_in_x_1_bits_wxd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_1_bits_reg_idxw = io_in_x_1_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_1_bits_warp_id = io_in_x_1_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_2_valid = io_in_x_2_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_x_io_in_2_bits_wb_wxd_rd = io_in_x_2_bits_wb_wxd_rd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_2_bits_wxd = io_in_x_2_bits_wxd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_2_bits_reg_idxw = io_in_x_2_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_2_bits_warp_id = io_in_x_2_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_3_valid = io_in_x_3_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_x_io_in_3_bits_wb_wxd_rd = io_in_x_3_bits_wb_wxd_rd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_3_bits_wxd = io_in_x_3_bits_wxd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_3_bits_reg_idxw = io_in_x_3_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_3_bits_warp_id = io_in_x_3_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_4_valid = io_in_x_4_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_x_io_in_4_bits_wb_wxd_rd = io_in_x_4_bits_wb_wxd_rd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_4_bits_wxd = io_in_x_4_bits_wxd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_4_bits_reg_idxw = io_in_x_4_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_x_io_in_4_bits_warp_id = io_in_x_4_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_valid = io_in_v_0_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_0 = io_in_v_0_bits_wb_wfd_rd_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_1 = io_in_v_0_bits_wb_wfd_rd_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_2 = io_in_v_0_bits_wb_wfd_rd_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_3 = io_in_v_0_bits_wb_wfd_rd_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_4 = io_in_v_0_bits_wb_wfd_rd_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_5 = io_in_v_0_bits_wb_wfd_rd_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_6 = io_in_v_0_bits_wb_wfd_rd_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wb_wfd_rd_7 = io_in_v_0_bits_wb_wfd_rd_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_0 = io_in_v_0_bits_wfd_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_1 = io_in_v_0_bits_wfd_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_2 = io_in_v_0_bits_wfd_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_3 = io_in_v_0_bits_wfd_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_4 = io_in_v_0_bits_wfd_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_5 = io_in_v_0_bits_wfd_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_6 = io_in_v_0_bits_wfd_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd_mask_7 = io_in_v_0_bits_wfd_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_wfd = io_in_v_0_bits_wfd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_reg_idxw = io_in_v_0_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_0_bits_warp_id = io_in_v_0_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_valid = io_in_v_1_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_0 = io_in_v_1_bits_wb_wfd_rd_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_1 = io_in_v_1_bits_wb_wfd_rd_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_2 = io_in_v_1_bits_wb_wfd_rd_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_3 = io_in_v_1_bits_wb_wfd_rd_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_4 = io_in_v_1_bits_wb_wfd_rd_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_5 = io_in_v_1_bits_wb_wfd_rd_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_6 = io_in_v_1_bits_wb_wfd_rd_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wb_wfd_rd_7 = io_in_v_1_bits_wb_wfd_rd_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_0 = io_in_v_1_bits_wfd_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_1 = io_in_v_1_bits_wfd_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_2 = io_in_v_1_bits_wfd_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_3 = io_in_v_1_bits_wfd_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_4 = io_in_v_1_bits_wfd_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_5 = io_in_v_1_bits_wfd_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_6 = io_in_v_1_bits_wfd_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd_mask_7 = io_in_v_1_bits_wfd_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_wfd = io_in_v_1_bits_wfd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_reg_idxw = io_in_v_1_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_1_bits_warp_id = io_in_v_1_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_valid = io_in_v_2_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_0 = io_in_v_2_bits_wb_wfd_rd_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_1 = io_in_v_2_bits_wb_wfd_rd_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_2 = io_in_v_2_bits_wb_wfd_rd_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_3 = io_in_v_2_bits_wb_wfd_rd_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_4 = io_in_v_2_bits_wb_wfd_rd_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_5 = io_in_v_2_bits_wb_wfd_rd_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_6 = io_in_v_2_bits_wb_wfd_rd_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wb_wfd_rd_7 = io_in_v_2_bits_wb_wfd_rd_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_0 = io_in_v_2_bits_wfd_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_1 = io_in_v_2_bits_wfd_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_2 = io_in_v_2_bits_wfd_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_3 = io_in_v_2_bits_wfd_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_4 = io_in_v_2_bits_wfd_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_5 = io_in_v_2_bits_wfd_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_6 = io_in_v_2_bits_wfd_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd_mask_7 = io_in_v_2_bits_wfd_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_wfd = io_in_v_2_bits_wfd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_reg_idxw = io_in_v_2_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_2_bits_warp_id = io_in_v_2_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_valid = io_in_v_3_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_0 = io_in_v_3_bits_wb_wfd_rd_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_1 = io_in_v_3_bits_wb_wfd_rd_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_2 = io_in_v_3_bits_wb_wfd_rd_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_3 = io_in_v_3_bits_wb_wfd_rd_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_4 = io_in_v_3_bits_wb_wfd_rd_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_5 = io_in_v_3_bits_wb_wfd_rd_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_6 = io_in_v_3_bits_wb_wfd_rd_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wb_wfd_rd_7 = io_in_v_3_bits_wb_wfd_rd_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_0 = io_in_v_3_bits_wfd_mask_0; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_1 = io_in_v_3_bits_wfd_mask_1; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_2 = io_in_v_3_bits_wfd_mask_2; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_3 = io_in_v_3_bits_wfd_mask_3; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_4 = io_in_v_3_bits_wfd_mask_4; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_5 = io_in_v_3_bits_wfd_mask_5; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_6 = io_in_v_3_bits_wfd_mask_6; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd_mask_7 = io_in_v_3_bits_wfd_mask_7; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_wfd = io_in_v_3_bits_wfd; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_reg_idxw = io_in_v_3_bits_reg_idxw; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_v_io_in_3_bits_warp_id = io_in_v_3_bits_warp_id; // @[Decoupled.scala 355:21 357:16]
endmodule
module Scoreboard(
  input        clock,
  input        reset,
  input  [1:0] io_ibuffer_if_ctrl_sel_alu2,
  input  [1:0] io_ibuffer_if_ctrl_sel_alu1,
  input        io_ibuffer_if_ctrl_isvec,
  input  [1:0] io_ibuffer_if_ctrl_sel_alu3,
  input        io_ibuffer_if_ctrl_mask,
  input        io_ibuffer_if_ctrl_mem,
  input  [4:0] io_ibuffer_if_ctrl_reg_idx1,
  input  [4:0] io_ibuffer_if_ctrl_reg_idx2,
  input  [4:0] io_ibuffer_if_ctrl_reg_idx3,
  input  [1:0] io_if_ctrl_branch,
  input        io_if_ctrl_barrier,
  input  [4:0] io_if_ctrl_reg_idxw,
  input        io_if_ctrl_wfd,
  input        io_if_ctrl_fence,
  input        io_if_ctrl_wxd,
  input        io_wb_v_ctrl_wfd,
  input  [4:0] io_wb_v_ctrl_reg_idxw,
  input        io_wb_x_ctrl_wxd,
  input  [4:0] io_wb_x_ctrl_reg_idxw,
  input        io_if_fire,
  input        io_br_ctrl,
  input        io_fence_end,
  input        io_wb_v_fire,
  input        io_wb_x_fire,
  output       io_delay
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] _r; // @[scoreboard.scala 69:27]
  reg [31:0] _r_1; // @[scoreboard.scala 69:27]
  wire [31:0] r = {_r_1[31:1], 1'h0}; // @[scoreboard.scala 70:37]
  reg  readb; // @[scoreboard.scala 69:27]
  reg  _r_3; // @[scoreboard.scala 69:27]
  wire  _T = io_if_fire & io_if_ctrl_wfd; // @[scoreboard.scala 86:28]
  wire [31:0] _T_1 = 32'h1 << io_if_ctrl_reg_idxw; // @[scoreboard.scala 73:57]
  wire [31:0] _T_2 = _T ? _T_1 : 32'h0; // @[scoreboard.scala 73:47]
  wire [31:0] _T_3 = _r | _T_2; // @[scoreboard.scala 65:67]
  wire  _T_5 = io_wb_v_fire & io_wb_v_ctrl_wfd; // @[scoreboard.scala 87:32]
  wire [31:0] _T_6 = 32'h1 << io_wb_v_ctrl_reg_idxw; // @[scoreboard.scala 73:57]
  wire [31:0] _T_7 = _T_5 ? _T_6 : 32'h0; // @[scoreboard.scala 73:47]
  wire [31:0] _T_8 = ~_T_7; // @[scoreboard.scala 66:72]
  wire [31:0] _T_9 = _T_3 & _T_8; // @[scoreboard.scala 66:69]
  wire  _T_10 = _T | _T_5; // @[scoreboard.scala 76:15]
  wire  _T_11 = io_if_fire & io_if_ctrl_wxd; // @[scoreboard.scala 88:28]
  wire [31:0] _T_13 = _T_11 ? _T_1 : 32'h0; // @[scoreboard.scala 73:47]
  wire [31:0] _T_14 = r | _T_13; // @[scoreboard.scala 65:67]
  wire  _T_16 = io_wb_x_fire & io_wb_x_ctrl_wxd; // @[scoreboard.scala 89:32]
  wire [31:0] _T_17 = 32'h1 << io_wb_x_ctrl_reg_idxw; // @[scoreboard.scala 73:57]
  wire [31:0] _T_18 = _T_16 ? _T_17 : 32'h0; // @[scoreboard.scala 73:47]
  wire [31:0] _T_19 = ~_T_18; // @[scoreboard.scala 66:72]
  wire [31:0] _T_20 = _T_14 & _T_19; // @[scoreboard.scala 66:69]
  wire  _T_21 = _T_11 | _T_16; // @[scoreboard.scala 76:15]
  wire  _T_24 = io_if_fire & (io_if_ctrl_branch != 2'h0 | io_if_ctrl_barrier); // @[scoreboard.scala 90:25]
  wire [1:0] _T_26 = _T_24 ? 2'h1 : 2'h0; // @[scoreboard.scala 73:47]
  wire [1:0] _GEN_8 = {{1'd0}, readb}; // @[scoreboard.scala 65:67]
  wire [1:0] _T_27 = _GEN_8 | _T_26; // @[scoreboard.scala 65:67]
  wire [1:0] _GEN_4 = _T_24 ? _T_27 : {{1'd0}, readb}; // @[scoreboard.scala 77:{16,21} 69:27]
  wire [1:0] _T_30 = io_br_ctrl ? 2'h1 : 2'h0; // @[scoreboard.scala 73:47]
  wire [1:0] _T_31 = ~_T_30; // @[scoreboard.scala 66:72]
  wire [1:0] _T_32 = _T_27 & _T_31; // @[scoreboard.scala 66:69]
  wire  _T_33 = _T_24 | io_br_ctrl; // @[scoreboard.scala 76:15]
  wire [1:0] _GEN_5 = _T_33 ? _T_32 : _GEN_4; // @[scoreboard.scala 77:{16,21}]
  wire  _T_34 = io_if_fire & io_if_ctrl_fence; // @[scoreboard.scala 92:27]
  wire [1:0] _T_36 = _T_34 ? 2'h1 : 2'h0; // @[scoreboard.scala 73:47]
  wire [1:0] _GEN_9 = {{1'd0}, _r_3}; // @[scoreboard.scala 65:67]
  wire [1:0] _T_37 = _GEN_9 | _T_36; // @[scoreboard.scala 65:67]
  wire [1:0] _GEN_6 = _T_34 ? _T_37 : {{1'd0}, _r_3}; // @[scoreboard.scala 77:{16,21} 69:27]
  wire [1:0] _T_40 = io_fence_end ? 2'h1 : 2'h0; // @[scoreboard.scala 73:47]
  wire [1:0] _T_41 = ~_T_40; // @[scoreboard.scala 66:72]
  wire [1:0] _T_42 = _T_37 & _T_41; // @[scoreboard.scala 66:69]
  wire  _T_43 = _T_34 | io_fence_end; // @[scoreboard.scala 76:15]
  wire [1:0] _GEN_7 = _T_43 ? _T_42 : _GEN_6; // @[scoreboard.scala 77:{16,21}]
  wire [31:0] _read1_T = r >> io_ibuffer_if_ctrl_reg_idx1; // @[scoreboard.scala 67:33]
  wire [31:0] _read1_T_2 = _r >> io_ibuffer_if_ctrl_reg_idx1; // @[scoreboard.scala 67:33]
  wire  read1 = 2'h2 == io_ibuffer_if_ctrl_sel_alu1 ? _read1_T_2[0] : 2'h1 == io_ibuffer_if_ctrl_sel_alu1 & _read1_T[0]; // @[Mux.scala 81:58]
  wire [31:0] _read2_T = r >> io_ibuffer_if_ctrl_reg_idx2; // @[scoreboard.scala 67:33]
  wire [31:0] _read2_T_2 = _r >> io_ibuffer_if_ctrl_reg_idx2; // @[scoreboard.scala 67:33]
  wire  read2 = 2'h2 == io_ibuffer_if_ctrl_sel_alu2 ? _read2_T_2[0] : 2'h1 == io_ibuffer_if_ctrl_sel_alu2 & _read2_T[0]; // @[Mux.scala 81:58]
  wire [31:0] _read3_T = _r >> io_ibuffer_if_ctrl_reg_idx3; // @[scoreboard.scala 67:33]
  wire  _read3_T_6 = io_ibuffer_if_ctrl_isvec ? _read3_T[0] : _read2_T[0]; // @[scoreboard.scala 96:128]
  wire  read3 = 2'h3 == io_ibuffer_if_ctrl_sel_alu3 ? _read3_T_6 : 2'h1 == io_ibuffer_if_ctrl_sel_alu3 & _read3_T[0]; // @[Mux.scala 81:58]
  wire  readm = io_ibuffer_if_ctrl_mask & _r[0]; // @[scoreboard.scala 97:16]
  wire  readf = io_ibuffer_if_ctrl_mem & _r_3; // @[scoreboard.scala 100:36]
  wire [1:0] _GEN_10 = reset ? 2'h0 : _GEN_5; // @[scoreboard.scala 69:{27,27}]
  wire [1:0] _GEN_11 = reset ? 2'h0 : _GEN_7; // @[scoreboard.scala 69:{27,27}]
  assign io_delay = read1 | read2 | read3 | readm | readb | readf; // @[scoreboard.scala 101:42]
  always @(posedge clock) begin
    if (reset) begin // @[scoreboard.scala 69:27]
      _r <= 32'h0; // @[scoreboard.scala 69:27]
    end else if (_T_10) begin // @[scoreboard.scala 77:16]
      _r <= _T_9; // @[scoreboard.scala 77:21]
    end else if (_T) begin // @[scoreboard.scala 77:16]
      _r <= _T_3; // @[scoreboard.scala 77:21]
    end
    if (reset) begin // @[scoreboard.scala 69:27]
      _r_1 <= 32'h0; // @[scoreboard.scala 69:27]
    end else if (_T_21) begin // @[scoreboard.scala 77:16]
      _r_1 <= _T_20; // @[scoreboard.scala 77:21]
    end else if (_T_11) begin // @[scoreboard.scala 77:16]
      _r_1 <= _T_14; // @[scoreboard.scala 77:21]
    end
    readb <= _GEN_10[0]; // @[scoreboard.scala 69:{27,27}]
    _r_3 <= _GEN_11[0]; // @[scoreboard.scala 69:{27,27}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _r = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _r_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  readb = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _r_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueWithFlush(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_inst,
  input  [1:0]  io_enq_bits_wid,
  input         io_enq_bits_fp,
  input  [1:0]  io_enq_bits_branch,
  input         io_enq_bits_simt_stack,
  input         io_enq_bits_simt_stack_op,
  input         io_enq_bits_barrier,
  input  [1:0]  io_enq_bits_csr,
  input         io_enq_bits_reverse,
  input  [1:0]  io_enq_bits_sel_alu2,
  input  [1:0]  io_enq_bits_sel_alu1,
  input         io_enq_bits_isvec,
  input  [1:0]  io_enq_bits_sel_alu3,
  input         io_enq_bits_mask,
  input  [2:0]  io_enq_bits_sel_imm,
  input         io_enq_bits_mem_unsigned,
  input  [5:0]  io_enq_bits_alu_fn,
  input         io_enq_bits_mem,
  input  [1:0]  io_enq_bits_mem_cmd,
  input  [1:0]  io_enq_bits_mop,
  input  [4:0]  io_enq_bits_reg_idx1,
  input  [4:0]  io_enq_bits_reg_idx2,
  input  [4:0]  io_enq_bits_reg_idx3,
  input  [4:0]  io_enq_bits_reg_idxw,
  input         io_enq_bits_wfd,
  input         io_enq_bits_fence,
  input         io_enq_bits_sfu,
  input         io_enq_bits_readmask,
  input         io_enq_bits_writemask,
  input         io_enq_bits_wxd,
  input  [31:0] io_enq_bits_pc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_inst,
  output [1:0]  io_deq_bits_wid,
  output        io_deq_bits_fp,
  output [1:0]  io_deq_bits_branch,
  output        io_deq_bits_simt_stack,
  output        io_deq_bits_simt_stack_op,
  output        io_deq_bits_barrier,
  output [1:0]  io_deq_bits_csr,
  output        io_deq_bits_reverse,
  output [1:0]  io_deq_bits_sel_alu2,
  output [1:0]  io_deq_bits_sel_alu1,
  output        io_deq_bits_isvec,
  output [1:0]  io_deq_bits_sel_alu3,
  output        io_deq_bits_mask,
  output [2:0]  io_deq_bits_sel_imm,
  output        io_deq_bits_mem_unsigned,
  output [5:0]  io_deq_bits_alu_fn,
  output        io_deq_bits_mem,
  output [1:0]  io_deq_bits_mem_cmd,
  output [1:0]  io_deq_bits_mop,
  output [4:0]  io_deq_bits_reg_idx1,
  output [4:0]  io_deq_bits_reg_idx2,
  output [4:0]  io_deq_bits_reg_idx3,
  output [4:0]  io_deq_bits_reg_idxw,
  output        io_deq_bits_wfd,
  output        io_deq_bits_fence,
  output        io_deq_bits_sfu,
  output        io_deq_bits_readmask,
  output        io_deq_bits_writemask,
  output        io_deq_bits_wxd,
  output [31:0] io_deq_bits_pc,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_inst [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_inst_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_inst_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [31:0] ram_inst_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [31:0] ram_inst_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_inst_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_inst_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_inst_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_wid [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_wid_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_wid_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_wid_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_wid_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_wid_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_wid_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_wid_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_fp [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_fp_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_branch [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_branch_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_branch_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_branch_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_branch_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_branch_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_branch_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_branch_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_simt_stack [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_simt_stack_op [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_simt_stack_op_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_barrier [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_barrier_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_csr [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_csr_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_csr_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_csr_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_csr_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_csr_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_csr_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_csr_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_reverse [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_reverse_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_sel_alu2 [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu2_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu2_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_sel_alu2_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_sel_alu2_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu2_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu2_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu2_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_sel_alu1 [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu1_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu1_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_sel_alu1_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_sel_alu1_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu1_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu1_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu1_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_isvec [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_isvec_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_sel_alu3 [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu3_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu3_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_sel_alu3_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_sel_alu3_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu3_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu3_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_alu3_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_mask [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_mask_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [2:0] ram_sel_imm [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_imm_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_imm_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [2:0] ram_sel_imm_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [2:0] ram_sel_imm_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_imm_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_imm_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_sel_imm_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_mem_unsigned [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_unsigned_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [5:0] ram_alu_fn [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_alu_fn_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_alu_fn_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [5:0] ram_alu_fn_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [5:0] ram_alu_fn_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_alu_fn_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_alu_fn_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_alu_fn_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_mem [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_mem_cmd [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_cmd_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_cmd_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_mem_cmd_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_mem_cmd_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_cmd_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_cmd_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_mem_cmd_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [1:0] ram_mop [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_mop_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_mop_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_mop_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [1:0] ram_mop_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_mop_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_mop_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_mop_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [4:0] ram_reg_idx1 [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx1_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx1_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idx1_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idx1_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx1_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx1_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx1_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [4:0] ram_reg_idx2 [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx2_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx2_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idx2_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idx2_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx2_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx2_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx2_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [4:0] ram_reg_idx3 [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx3_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx3_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idx3_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idx3_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx3_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx3_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idx3_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [4:0] ram_reg_idxw [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idxw_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idxw_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idxw_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [4:0] ram_reg_idxw_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idxw_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idxw_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_reg_idxw_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_wfd [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_wfd_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_fence [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_fence_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_sfu [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_sfu_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_readmask [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_readmask_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_writemask [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_writemask_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  ram_wxd [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_wxd_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg [31:0] ram_pc [0:1]; // @[QueueWithFlush.scala 303:95]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[QueueWithFlush.scala 303:95]
  wire  ram_pc_io_deq_bits_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire [31:0] ram_pc_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire [31:0] ram_pc_MPORT_data; // @[QueueWithFlush.scala 303:95]
  wire  ram_pc_MPORT_addr; // @[QueueWithFlush.scala 303:95]
  wire  ram_pc_MPORT_mask; // @[QueueWithFlush.scala 303:95]
  wire  ram_pc_MPORT_en; // @[QueueWithFlush.scala 303:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[QueueWithFlush.scala 306:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[QueueWithFlush.scala 307:33]
  wire  empty = ptr_match & ~maybe_full; // @[QueueWithFlush.scala 308:25]
  wire  full = ptr_match & maybe_full; // @[QueueWithFlush.scala 309:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_inst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_inst_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_inst_io_deq_bits_MPORT_data = ram_inst[ram_inst_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_inst_MPORT_data = io_enq_bits_inst;
  assign ram_inst_MPORT_addr = enq_ptr_value;
  assign ram_inst_MPORT_mask = 1'h1;
  assign ram_inst_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wid_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_wid_io_deq_bits_MPORT_data = ram_wid[ram_wid_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_wid_MPORT_data = io_enq_bits_wid;
  assign ram_wid_MPORT_addr = enq_ptr_value;
  assign ram_wid_MPORT_mask = 1'h1;
  assign ram_wid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_fp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_fp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_fp_io_deq_bits_MPORT_data = ram_fp[ram_fp_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_fp_MPORT_data = io_enq_bits_fp;
  assign ram_fp_MPORT_addr = enq_ptr_value;
  assign ram_fp_MPORT_mask = 1'h1;
  assign ram_fp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_branch_io_deq_bits_MPORT_en = 1'h1;
  assign ram_branch_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_branch_io_deq_bits_MPORT_data = ram_branch[ram_branch_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_branch_MPORT_data = io_enq_bits_branch;
  assign ram_branch_MPORT_addr = enq_ptr_value;
  assign ram_branch_MPORT_mask = 1'h1;
  assign ram_branch_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_simt_stack_io_deq_bits_MPORT_en = 1'h1;
  assign ram_simt_stack_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_simt_stack_io_deq_bits_MPORT_data = ram_simt_stack[ram_simt_stack_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_simt_stack_MPORT_data = io_enq_bits_simt_stack;
  assign ram_simt_stack_MPORT_addr = enq_ptr_value;
  assign ram_simt_stack_MPORT_mask = 1'h1;
  assign ram_simt_stack_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_simt_stack_op_io_deq_bits_MPORT_en = 1'h1;
  assign ram_simt_stack_op_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_simt_stack_op_io_deq_bits_MPORT_data = ram_simt_stack_op[ram_simt_stack_op_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_simt_stack_op_MPORT_data = io_enq_bits_simt_stack_op;
  assign ram_simt_stack_op_MPORT_addr = enq_ptr_value;
  assign ram_simt_stack_op_MPORT_mask = 1'h1;
  assign ram_simt_stack_op_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_barrier_io_deq_bits_MPORT_en = 1'h1;
  assign ram_barrier_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_barrier_io_deq_bits_MPORT_data = ram_barrier[ram_barrier_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_barrier_MPORT_data = io_enq_bits_barrier;
  assign ram_barrier_MPORT_addr = enq_ptr_value;
  assign ram_barrier_MPORT_mask = 1'h1;
  assign ram_barrier_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_csr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_csr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_csr_io_deq_bits_MPORT_data = ram_csr[ram_csr_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_csr_MPORT_data = io_enq_bits_csr;
  assign ram_csr_MPORT_addr = enq_ptr_value;
  assign ram_csr_MPORT_mask = 1'h1;
  assign ram_csr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reverse_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reverse_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_reverse_io_deq_bits_MPORT_data = ram_reverse[ram_reverse_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_reverse_MPORT_data = io_enq_bits_reverse;
  assign ram_reverse_MPORT_addr = enq_ptr_value;
  assign ram_reverse_MPORT_mask = 1'h1;
  assign ram_reverse_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sel_alu2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_alu2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sel_alu2_io_deq_bits_MPORT_data = ram_sel_alu2[ram_sel_alu2_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_sel_alu2_MPORT_data = io_enq_bits_sel_alu2;
  assign ram_sel_alu2_MPORT_addr = enq_ptr_value;
  assign ram_sel_alu2_MPORT_mask = 1'h1;
  assign ram_sel_alu2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sel_alu1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_alu1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sel_alu1_io_deq_bits_MPORT_data = ram_sel_alu1[ram_sel_alu1_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_sel_alu1_MPORT_data = io_enq_bits_sel_alu1;
  assign ram_sel_alu1_MPORT_addr = enq_ptr_value;
  assign ram_sel_alu1_MPORT_mask = 1'h1;
  assign ram_sel_alu1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_isvec_io_deq_bits_MPORT_en = 1'h1;
  assign ram_isvec_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_isvec_io_deq_bits_MPORT_data = ram_isvec[ram_isvec_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_isvec_MPORT_data = io_enq_bits_isvec;
  assign ram_isvec_MPORT_addr = enq_ptr_value;
  assign ram_isvec_MPORT_mask = 1'h1;
  assign ram_isvec_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sel_alu3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_alu3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sel_alu3_io_deq_bits_MPORT_data = ram_sel_alu3[ram_sel_alu3_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_sel_alu3_MPORT_data = io_enq_bits_sel_alu3;
  assign ram_sel_alu3_MPORT_addr = enq_ptr_value;
  assign ram_sel_alu3_MPORT_mask = 1'h1;
  assign ram_sel_alu3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sel_imm_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sel_imm_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sel_imm_io_deq_bits_MPORT_data = ram_sel_imm[ram_sel_imm_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_sel_imm_MPORT_data = io_enq_bits_sel_imm;
  assign ram_sel_imm_MPORT_addr = enq_ptr_value;
  assign ram_sel_imm_MPORT_mask = 1'h1;
  assign ram_sel_imm_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mem_unsigned_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mem_unsigned_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mem_unsigned_io_deq_bits_MPORT_data = ram_mem_unsigned[ram_mem_unsigned_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_mem_unsigned_MPORT_data = io_enq_bits_mem_unsigned;
  assign ram_mem_unsigned_MPORT_addr = enq_ptr_value;
  assign ram_mem_unsigned_MPORT_mask = 1'h1;
  assign ram_mem_unsigned_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_alu_fn_io_deq_bits_MPORT_en = 1'h1;
  assign ram_alu_fn_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_alu_fn_io_deq_bits_MPORT_data = ram_alu_fn[ram_alu_fn_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_alu_fn_MPORT_data = io_enq_bits_alu_fn;
  assign ram_alu_fn_MPORT_addr = enq_ptr_value;
  assign ram_alu_fn_MPORT_mask = 1'h1;
  assign ram_alu_fn_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mem_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mem_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mem_io_deq_bits_MPORT_data = ram_mem[ram_mem_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_mem_MPORT_data = io_enq_bits_mem;
  assign ram_mem_MPORT_addr = enq_ptr_value;
  assign ram_mem_MPORT_mask = 1'h1;
  assign ram_mem_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mem_cmd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mem_cmd_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mem_cmd_io_deq_bits_MPORT_data = ram_mem_cmd[ram_mem_cmd_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_mem_cmd_MPORT_data = io_enq_bits_mem_cmd;
  assign ram_mem_cmd_MPORT_addr = enq_ptr_value;
  assign ram_mem_cmd_MPORT_mask = 1'h1;
  assign ram_mem_cmd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mop_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mop_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mop_io_deq_bits_MPORT_data = ram_mop[ram_mop_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_mop_MPORT_data = io_enq_bits_mop;
  assign ram_mop_MPORT_addr = enq_ptr_value;
  assign ram_mop_MPORT_mask = 1'h1;
  assign ram_mop_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reg_idx1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reg_idx1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_reg_idx1_io_deq_bits_MPORT_data = ram_reg_idx1[ram_reg_idx1_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_reg_idx1_MPORT_data = io_enq_bits_reg_idx1;
  assign ram_reg_idx1_MPORT_addr = enq_ptr_value;
  assign ram_reg_idx1_MPORT_mask = 1'h1;
  assign ram_reg_idx1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reg_idx2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reg_idx2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_reg_idx2_io_deq_bits_MPORT_data = ram_reg_idx2[ram_reg_idx2_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_reg_idx2_MPORT_data = io_enq_bits_reg_idx2;
  assign ram_reg_idx2_MPORT_addr = enq_ptr_value;
  assign ram_reg_idx2_MPORT_mask = 1'h1;
  assign ram_reg_idx2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reg_idx3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reg_idx3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_reg_idx3_io_deq_bits_MPORT_data = ram_reg_idx3[ram_reg_idx3_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_reg_idx3_MPORT_data = io_enq_bits_reg_idx3;
  assign ram_reg_idx3_MPORT_addr = enq_ptr_value;
  assign ram_reg_idx3_MPORT_mask = 1'h1;
  assign ram_reg_idx3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_reg_idxw_io_deq_bits_MPORT_en = 1'h1;
  assign ram_reg_idxw_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_reg_idxw_io_deq_bits_MPORT_data = ram_reg_idxw[ram_reg_idxw_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_reg_idxw_MPORT_data = io_enq_bits_reg_idxw;
  assign ram_reg_idxw_MPORT_addr = enq_ptr_value;
  assign ram_reg_idxw_MPORT_mask = 1'h1;
  assign ram_reg_idxw_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wfd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wfd_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_wfd_io_deq_bits_MPORT_data = ram_wfd[ram_wfd_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_wfd_MPORT_data = io_enq_bits_wfd;
  assign ram_wfd_MPORT_addr = enq_ptr_value;
  assign ram_wfd_MPORT_mask = 1'h1;
  assign ram_wfd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_fence_io_deq_bits_MPORT_en = 1'h1;
  assign ram_fence_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_fence_io_deq_bits_MPORT_data = ram_fence[ram_fence_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_fence_MPORT_data = io_enq_bits_fence;
  assign ram_fence_MPORT_addr = enq_ptr_value;
  assign ram_fence_MPORT_mask = 1'h1;
  assign ram_fence_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sfu_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sfu_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sfu_io_deq_bits_MPORT_data = ram_sfu[ram_sfu_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_sfu_MPORT_data = io_enq_bits_sfu;
  assign ram_sfu_MPORT_addr = enq_ptr_value;
  assign ram_sfu_MPORT_mask = 1'h1;
  assign ram_sfu_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_readmask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_readmask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_readmask_io_deq_bits_MPORT_data = ram_readmask[ram_readmask_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_readmask_MPORT_data = io_enq_bits_readmask;
  assign ram_readmask_MPORT_addr = enq_ptr_value;
  assign ram_readmask_MPORT_mask = 1'h1;
  assign ram_readmask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_writemask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_writemask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_writemask_io_deq_bits_MPORT_data = ram_writemask[ram_writemask_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_writemask_MPORT_data = io_enq_bits_writemask;
  assign ram_writemask_MPORT_addr = enq_ptr_value;
  assign ram_writemask_MPORT_mask = 1'h1;
  assign ram_writemask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_wxd_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wxd_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_wxd_io_deq_bits_MPORT_data = ram_wxd[ram_wxd_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_wxd_MPORT_data = io_enq_bits_wxd;
  assign ram_wxd_MPORT_addr = enq_ptr_value;
  assign ram_wxd_MPORT_mask = 1'h1;
  assign ram_wxd_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[QueueWithFlush.scala 303:95]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[QueueWithFlush.scala 333:19]
  assign io_deq_valid = ~empty; // @[QueueWithFlush.scala 332:19]
  assign io_deq_bits_inst = ram_inst_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_wid = ram_wid_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_fp = ram_fp_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_branch = ram_branch_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_simt_stack = ram_simt_stack_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_simt_stack_op = ram_simt_stack_op_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_barrier = ram_barrier_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_csr = ram_csr_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_reverse = ram_reverse_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_sel_alu2 = ram_sel_alu2_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_sel_alu1 = ram_sel_alu1_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_isvec = ram_isvec_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_sel_alu3 = ram_sel_alu3_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_sel_imm = ram_sel_imm_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_mem_unsigned = ram_mem_unsigned_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_alu_fn = ram_alu_fn_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_mem = ram_mem_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_mem_cmd = ram_mem_cmd_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_mop = ram_mop_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_reg_idx1 = ram_reg_idx1_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_reg_idx2 = ram_reg_idx2_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_reg_idx3 = ram_reg_idx3_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_reg_idxw = ram_reg_idxw_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_wfd = ram_wfd_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_fence = ram_fence_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_sfu = ram_sfu_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_readmask = ram_readmask_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_writemask = ram_writemask_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_wxd = ram_wxd_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[QueueWithFlush.scala 340:17]
  always @(posedge clock) begin
    if (ram_inst_MPORT_en & ram_inst_MPORT_mask) begin
      ram_inst[ram_inst_MPORT_addr] <= ram_inst_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_wid_MPORT_en & ram_wid_MPORT_mask) begin
      ram_wid[ram_wid_MPORT_addr] <= ram_wid_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_fp_MPORT_en & ram_fp_MPORT_mask) begin
      ram_fp[ram_fp_MPORT_addr] <= ram_fp_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_branch_MPORT_en & ram_branch_MPORT_mask) begin
      ram_branch[ram_branch_MPORT_addr] <= ram_branch_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_simt_stack_MPORT_en & ram_simt_stack_MPORT_mask) begin
      ram_simt_stack[ram_simt_stack_MPORT_addr] <= ram_simt_stack_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_simt_stack_op_MPORT_en & ram_simt_stack_op_MPORT_mask) begin
      ram_simt_stack_op[ram_simt_stack_op_MPORT_addr] <= ram_simt_stack_op_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_barrier_MPORT_en & ram_barrier_MPORT_mask) begin
      ram_barrier[ram_barrier_MPORT_addr] <= ram_barrier_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_csr_MPORT_en & ram_csr_MPORT_mask) begin
      ram_csr[ram_csr_MPORT_addr] <= ram_csr_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_reverse_MPORT_en & ram_reverse_MPORT_mask) begin
      ram_reverse[ram_reverse_MPORT_addr] <= ram_reverse_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_sel_alu2_MPORT_en & ram_sel_alu2_MPORT_mask) begin
      ram_sel_alu2[ram_sel_alu2_MPORT_addr] <= ram_sel_alu2_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_sel_alu1_MPORT_en & ram_sel_alu1_MPORT_mask) begin
      ram_sel_alu1[ram_sel_alu1_MPORT_addr] <= ram_sel_alu1_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_isvec_MPORT_en & ram_isvec_MPORT_mask) begin
      ram_isvec[ram_isvec_MPORT_addr] <= ram_isvec_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_sel_alu3_MPORT_en & ram_sel_alu3_MPORT_mask) begin
      ram_sel_alu3[ram_sel_alu3_MPORT_addr] <= ram_sel_alu3_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_sel_imm_MPORT_en & ram_sel_imm_MPORT_mask) begin
      ram_sel_imm[ram_sel_imm_MPORT_addr] <= ram_sel_imm_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_mem_unsigned_MPORT_en & ram_mem_unsigned_MPORT_mask) begin
      ram_mem_unsigned[ram_mem_unsigned_MPORT_addr] <= ram_mem_unsigned_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_alu_fn_MPORT_en & ram_alu_fn_MPORT_mask) begin
      ram_alu_fn[ram_alu_fn_MPORT_addr] <= ram_alu_fn_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_mem_MPORT_en & ram_mem_MPORT_mask) begin
      ram_mem[ram_mem_MPORT_addr] <= ram_mem_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_mem_cmd_MPORT_en & ram_mem_cmd_MPORT_mask) begin
      ram_mem_cmd[ram_mem_cmd_MPORT_addr] <= ram_mem_cmd_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_mop_MPORT_en & ram_mop_MPORT_mask) begin
      ram_mop[ram_mop_MPORT_addr] <= ram_mop_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_reg_idx1_MPORT_en & ram_reg_idx1_MPORT_mask) begin
      ram_reg_idx1[ram_reg_idx1_MPORT_addr] <= ram_reg_idx1_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_reg_idx2_MPORT_en & ram_reg_idx2_MPORT_mask) begin
      ram_reg_idx2[ram_reg_idx2_MPORT_addr] <= ram_reg_idx2_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_reg_idx3_MPORT_en & ram_reg_idx3_MPORT_mask) begin
      ram_reg_idx3[ram_reg_idx3_MPORT_addr] <= ram_reg_idx3_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_reg_idxw_MPORT_en & ram_reg_idxw_MPORT_mask) begin
      ram_reg_idxw[ram_reg_idxw_MPORT_addr] <= ram_reg_idxw_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_wfd_MPORT_en & ram_wfd_MPORT_mask) begin
      ram_wfd[ram_wfd_MPORT_addr] <= ram_wfd_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_fence_MPORT_en & ram_fence_MPORT_mask) begin
      ram_fence[ram_fence_MPORT_addr] <= ram_fence_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_sfu_MPORT_en & ram_sfu_MPORT_mask) begin
      ram_sfu[ram_sfu_MPORT_addr] <= ram_sfu_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_readmask_MPORT_en & ram_readmask_MPORT_mask) begin
      ram_readmask[ram_readmask_MPORT_addr] <= ram_readmask_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_writemask_MPORT_en & ram_writemask_MPORT_mask) begin
      ram_writemask[ram_writemask_MPORT_addr] <= ram_writemask_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_wxd_MPORT_en & ram_wxd_MPORT_mask) begin
      ram_wxd[ram_wxd_MPORT_addr] <= ram_wxd_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[QueueWithFlush.scala 303:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_flush) begin // @[QueueWithFlush.scala 326:15]
      enq_ptr_value <= 1'h0; // @[Counter.scala 99:11]
    end else if (do_enq) begin // @[QueueWithFlush.scala 316:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_flush) begin // @[QueueWithFlush.scala 326:15]
      deq_ptr_value <= 1'h0; // @[Counter.scala 99:11]
    end else if (do_deq) begin // @[QueueWithFlush.scala 320:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[QueueWithFlush.scala 306:27]
      maybe_full <= 1'h0; // @[QueueWithFlush.scala 306:27]
    end else if (io_flush) begin // @[QueueWithFlush.scala 326:15]
      maybe_full <= 1'h0; // @[QueueWithFlush.scala 329:16]
    end else if (do_enq != do_deq) begin // @[QueueWithFlush.scala 323:27]
      maybe_full <= do_enq; // @[QueueWithFlush.scala 324:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_inst[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_wid[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_fp[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_branch[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_simt_stack[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_simt_stack_op[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_barrier[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_csr[initvar] = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_reverse[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sel_alu2[initvar] = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sel_alu1[initvar] = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_isvec[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sel_alu3[initvar] = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sel_imm[initvar] = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mem_unsigned[initvar] = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_alu_fn[initvar] = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mem[initvar] = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mem_cmd[initvar] = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mop[initvar] = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_reg_idx1[initvar] = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_reg_idx2[initvar] = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_reg_idx3[initvar] = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_reg_idxw[initvar] = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_wfd[initvar] = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_fence[initvar] = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sfu[initvar] = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_readmask[initvar] = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_writemask[initvar] = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_wxd[initvar] = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_pc[initvar] = _RAND_30[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  enq_ptr_value = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  deq_ptr_value = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  maybe_full = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module instbuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_inst,
  input  [1:0]  io_in_bits_wid,
  input         io_in_bits_fp,
  input  [1:0]  io_in_bits_branch,
  input         io_in_bits_simt_stack,
  input         io_in_bits_simt_stack_op,
  input         io_in_bits_barrier,
  input  [1:0]  io_in_bits_csr,
  input         io_in_bits_reverse,
  input  [1:0]  io_in_bits_sel_alu2,
  input  [1:0]  io_in_bits_sel_alu1,
  input         io_in_bits_isvec,
  input  [1:0]  io_in_bits_sel_alu3,
  input         io_in_bits_mask,
  input  [2:0]  io_in_bits_sel_imm,
  input         io_in_bits_mem_unsigned,
  input  [5:0]  io_in_bits_alu_fn,
  input         io_in_bits_mem,
  input  [1:0]  io_in_bits_mem_cmd,
  input  [1:0]  io_in_bits_mop,
  input  [4:0]  io_in_bits_reg_idx1,
  input  [4:0]  io_in_bits_reg_idx2,
  input  [4:0]  io_in_bits_reg_idx3,
  input  [4:0]  io_in_bits_reg_idxw,
  input         io_in_bits_wfd,
  input         io_in_bits_fence,
  input         io_in_bits_sfu,
  input         io_in_bits_readmask,
  input         io_in_bits_writemask,
  input         io_in_bits_wxd,
  input  [31:0] io_in_bits_pc,
  input         io_flush_valid,
  input  [1:0]  io_flush_bits,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [31:0] io_out_0_bits_inst,
  output [1:0]  io_out_0_bits_wid,
  output        io_out_0_bits_fp,
  output [1:0]  io_out_0_bits_branch,
  output        io_out_0_bits_simt_stack,
  output        io_out_0_bits_simt_stack_op,
  output        io_out_0_bits_barrier,
  output [1:0]  io_out_0_bits_csr,
  output        io_out_0_bits_reverse,
  output [1:0]  io_out_0_bits_sel_alu2,
  output [1:0]  io_out_0_bits_sel_alu1,
  output        io_out_0_bits_isvec,
  output [1:0]  io_out_0_bits_sel_alu3,
  output        io_out_0_bits_mask,
  output [2:0]  io_out_0_bits_sel_imm,
  output        io_out_0_bits_mem_unsigned,
  output [5:0]  io_out_0_bits_alu_fn,
  output        io_out_0_bits_mem,
  output [1:0]  io_out_0_bits_mem_cmd,
  output [1:0]  io_out_0_bits_mop,
  output [4:0]  io_out_0_bits_reg_idx1,
  output [4:0]  io_out_0_bits_reg_idx2,
  output [4:0]  io_out_0_bits_reg_idx3,
  output [4:0]  io_out_0_bits_reg_idxw,
  output        io_out_0_bits_wfd,
  output        io_out_0_bits_fence,
  output        io_out_0_bits_sfu,
  output        io_out_0_bits_readmask,
  output        io_out_0_bits_writemask,
  output        io_out_0_bits_wxd,
  output [31:0] io_out_0_bits_pc,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [31:0] io_out_1_bits_inst,
  output [1:0]  io_out_1_bits_wid,
  output        io_out_1_bits_fp,
  output [1:0]  io_out_1_bits_branch,
  output        io_out_1_bits_simt_stack,
  output        io_out_1_bits_simt_stack_op,
  output        io_out_1_bits_barrier,
  output [1:0]  io_out_1_bits_csr,
  output        io_out_1_bits_reverse,
  output [1:0]  io_out_1_bits_sel_alu2,
  output [1:0]  io_out_1_bits_sel_alu1,
  output        io_out_1_bits_isvec,
  output [1:0]  io_out_1_bits_sel_alu3,
  output        io_out_1_bits_mask,
  output [2:0]  io_out_1_bits_sel_imm,
  output        io_out_1_bits_mem_unsigned,
  output [5:0]  io_out_1_bits_alu_fn,
  output        io_out_1_bits_mem,
  output [1:0]  io_out_1_bits_mem_cmd,
  output [1:0]  io_out_1_bits_mop,
  output [4:0]  io_out_1_bits_reg_idx1,
  output [4:0]  io_out_1_bits_reg_idx2,
  output [4:0]  io_out_1_bits_reg_idx3,
  output [4:0]  io_out_1_bits_reg_idxw,
  output        io_out_1_bits_wfd,
  output        io_out_1_bits_fence,
  output        io_out_1_bits_sfu,
  output        io_out_1_bits_readmask,
  output        io_out_1_bits_writemask,
  output        io_out_1_bits_wxd,
  output [31:0] io_out_1_bits_pc,
  input         io_out_2_ready,
  output        io_out_2_valid,
  output [31:0] io_out_2_bits_inst,
  output [1:0]  io_out_2_bits_wid,
  output        io_out_2_bits_fp,
  output [1:0]  io_out_2_bits_branch,
  output        io_out_2_bits_simt_stack,
  output        io_out_2_bits_simt_stack_op,
  output        io_out_2_bits_barrier,
  output [1:0]  io_out_2_bits_csr,
  output        io_out_2_bits_reverse,
  output [1:0]  io_out_2_bits_sel_alu2,
  output [1:0]  io_out_2_bits_sel_alu1,
  output        io_out_2_bits_isvec,
  output [1:0]  io_out_2_bits_sel_alu3,
  output        io_out_2_bits_mask,
  output [2:0]  io_out_2_bits_sel_imm,
  output        io_out_2_bits_mem_unsigned,
  output [5:0]  io_out_2_bits_alu_fn,
  output        io_out_2_bits_mem,
  output [1:0]  io_out_2_bits_mem_cmd,
  output [1:0]  io_out_2_bits_mop,
  output [4:0]  io_out_2_bits_reg_idx1,
  output [4:0]  io_out_2_bits_reg_idx2,
  output [4:0]  io_out_2_bits_reg_idx3,
  output [4:0]  io_out_2_bits_reg_idxw,
  output        io_out_2_bits_wfd,
  output        io_out_2_bits_fence,
  output        io_out_2_bits_sfu,
  output        io_out_2_bits_readmask,
  output        io_out_2_bits_writemask,
  output        io_out_2_bits_wxd,
  output [31:0] io_out_2_bits_pc,
  input         io_out_3_ready,
  output        io_out_3_valid,
  output [31:0] io_out_3_bits_inst,
  output [1:0]  io_out_3_bits_wid,
  output        io_out_3_bits_fp,
  output [1:0]  io_out_3_bits_branch,
  output        io_out_3_bits_simt_stack,
  output        io_out_3_bits_simt_stack_op,
  output        io_out_3_bits_barrier,
  output [1:0]  io_out_3_bits_csr,
  output        io_out_3_bits_reverse,
  output [1:0]  io_out_3_bits_sel_alu2,
  output [1:0]  io_out_3_bits_sel_alu1,
  output        io_out_3_bits_isvec,
  output [1:0]  io_out_3_bits_sel_alu3,
  output        io_out_3_bits_mask,
  output [2:0]  io_out_3_bits_sel_imm,
  output        io_out_3_bits_mem_unsigned,
  output [5:0]  io_out_3_bits_alu_fn,
  output        io_out_3_bits_mem,
  output [1:0]  io_out_3_bits_mem_cmd,
  output [1:0]  io_out_3_bits_mop,
  output [4:0]  io_out_3_bits_reg_idx1,
  output [4:0]  io_out_3_bits_reg_idx2,
  output [4:0]  io_out_3_bits_reg_idx3,
  output [4:0]  io_out_3_bits_reg_idxw,
  output        io_out_3_bits_wfd,
  output        io_out_3_bits_fence,
  output        io_out_3_bits_sfu,
  output        io_out_3_bits_readmask,
  output        io_out_3_bits_writemask,
  output        io_out_3_bits_wxd,
  output [31:0] io_out_3_bits_pc,
  output        io_ibuffer_ready_0,
  output        io_ibuffer_ready_1,
  output        io_ibuffer_ready_2,
  output        io_ibuffer_ready_3
);
  wire  fifo_0_clock; // @[ibuffer.scala 20:24]
  wire  fifo_0_reset; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_0_io_enq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_0_io_enq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_0_io_enq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_enq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_enq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_enq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_enq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_enq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_enq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_0_io_enq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_0_io_deq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_0_io_deq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_0_io_deq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_0_io_deq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_deq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_deq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_deq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_0_io_deq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_deq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_0_io_deq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_0_io_flush; // @[ibuffer.scala 20:24]
  wire  fifo_1_clock; // @[ibuffer.scala 20:24]
  wire  fifo_1_reset; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_1_io_enq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_1_io_enq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_1_io_enq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_enq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_enq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_enq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_enq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_enq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_enq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_1_io_enq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_1_io_deq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_1_io_deq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_1_io_deq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_1_io_deq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_deq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_deq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_deq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_1_io_deq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_deq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_1_io_deq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_1_io_flush; // @[ibuffer.scala 20:24]
  wire  fifo_2_clock; // @[ibuffer.scala 20:24]
  wire  fifo_2_reset; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_2_io_enq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_2_io_enq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_2_io_enq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_enq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_enq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_enq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_enq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_enq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_enq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_2_io_enq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_2_io_deq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_2_io_deq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_2_io_deq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_2_io_deq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_deq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_deq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_deq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_2_io_deq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_deq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_2_io_deq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_2_io_flush; // @[ibuffer.scala 20:24]
  wire  fifo_3_clock; // @[ibuffer.scala 20:24]
  wire  fifo_3_reset; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_3_io_enq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_3_io_enq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_3_io_enq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_enq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_enq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_enq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_enq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_enq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_enq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_3_io_enq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_ready; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_valid; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_3_io_deq_bits_inst; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_wid; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_fp; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_branch; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_simt_stack; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_simt_stack_op; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_barrier; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_csr; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_reverse; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_sel_alu2; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_sel_alu1; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_isvec; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_sel_alu3; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_mask; // @[ibuffer.scala 20:24]
  wire [2:0] fifo_3_io_deq_bits_sel_imm; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_mem_unsigned; // @[ibuffer.scala 20:24]
  wire [5:0] fifo_3_io_deq_bits_alu_fn; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_mem; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_mem_cmd; // @[ibuffer.scala 20:24]
  wire [1:0] fifo_3_io_deq_bits_mop; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_deq_bits_reg_idx1; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_deq_bits_reg_idx2; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_deq_bits_reg_idx3; // @[ibuffer.scala 20:24]
  wire [4:0] fifo_3_io_deq_bits_reg_idxw; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_wfd; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_fence; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_sfu; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_readmask; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_writemask; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_deq_bits_wxd; // @[ibuffer.scala 20:24]
  wire [31:0] fifo_3_io_deq_bits_pc; // @[ibuffer.scala 20:24]
  wire  fifo_3_io_flush; // @[ibuffer.scala 20:24]
  wire  _x_single_io_enq_valid_T = 2'h0 == io_in_bits_wid; // @[ibuffer.scala 23:45]
  wire  _GEN_0 = _x_single_io_enq_valid_T & fifo_0_io_enq_ready; // @[ibuffer.scala 18:14 24:{40,52}]
  wire  _x_single_io_enq_valid_T_2 = 2'h1 == io_in_bits_wid; // @[ibuffer.scala 23:45]
  wire  _GEN_1 = _x_single_io_enq_valid_T_2 ? fifo_1_io_enq_ready : _GEN_0; // @[ibuffer.scala 24:{40,52}]
  wire  _x_single_io_enq_valid_T_4 = 2'h2 == io_in_bits_wid; // @[ibuffer.scala 23:45]
  wire  _GEN_2 = _x_single_io_enq_valid_T_4 ? fifo_2_io_enq_ready : _GEN_1; // @[ibuffer.scala 24:{40,52}]
  wire  _x_single_io_enq_valid_T_6 = 2'h3 == io_in_bits_wid; // @[ibuffer.scala 23:45]
  QueueWithFlush fifo_0 ( // @[ibuffer.scala 20:24]
    .clock(fifo_0_clock),
    .reset(fifo_0_reset),
    .io_enq_ready(fifo_0_io_enq_ready),
    .io_enq_valid(fifo_0_io_enq_valid),
    .io_enq_bits_inst(fifo_0_io_enq_bits_inst),
    .io_enq_bits_wid(fifo_0_io_enq_bits_wid),
    .io_enq_bits_fp(fifo_0_io_enq_bits_fp),
    .io_enq_bits_branch(fifo_0_io_enq_bits_branch),
    .io_enq_bits_simt_stack(fifo_0_io_enq_bits_simt_stack),
    .io_enq_bits_simt_stack_op(fifo_0_io_enq_bits_simt_stack_op),
    .io_enq_bits_barrier(fifo_0_io_enq_bits_barrier),
    .io_enq_bits_csr(fifo_0_io_enq_bits_csr),
    .io_enq_bits_reverse(fifo_0_io_enq_bits_reverse),
    .io_enq_bits_sel_alu2(fifo_0_io_enq_bits_sel_alu2),
    .io_enq_bits_sel_alu1(fifo_0_io_enq_bits_sel_alu1),
    .io_enq_bits_isvec(fifo_0_io_enq_bits_isvec),
    .io_enq_bits_sel_alu3(fifo_0_io_enq_bits_sel_alu3),
    .io_enq_bits_mask(fifo_0_io_enq_bits_mask),
    .io_enq_bits_sel_imm(fifo_0_io_enq_bits_sel_imm),
    .io_enq_bits_mem_unsigned(fifo_0_io_enq_bits_mem_unsigned),
    .io_enq_bits_alu_fn(fifo_0_io_enq_bits_alu_fn),
    .io_enq_bits_mem(fifo_0_io_enq_bits_mem),
    .io_enq_bits_mem_cmd(fifo_0_io_enq_bits_mem_cmd),
    .io_enq_bits_mop(fifo_0_io_enq_bits_mop),
    .io_enq_bits_reg_idx1(fifo_0_io_enq_bits_reg_idx1),
    .io_enq_bits_reg_idx2(fifo_0_io_enq_bits_reg_idx2),
    .io_enq_bits_reg_idx3(fifo_0_io_enq_bits_reg_idx3),
    .io_enq_bits_reg_idxw(fifo_0_io_enq_bits_reg_idxw),
    .io_enq_bits_wfd(fifo_0_io_enq_bits_wfd),
    .io_enq_bits_fence(fifo_0_io_enq_bits_fence),
    .io_enq_bits_sfu(fifo_0_io_enq_bits_sfu),
    .io_enq_bits_readmask(fifo_0_io_enq_bits_readmask),
    .io_enq_bits_writemask(fifo_0_io_enq_bits_writemask),
    .io_enq_bits_wxd(fifo_0_io_enq_bits_wxd),
    .io_enq_bits_pc(fifo_0_io_enq_bits_pc),
    .io_deq_ready(fifo_0_io_deq_ready),
    .io_deq_valid(fifo_0_io_deq_valid),
    .io_deq_bits_inst(fifo_0_io_deq_bits_inst),
    .io_deq_bits_wid(fifo_0_io_deq_bits_wid),
    .io_deq_bits_fp(fifo_0_io_deq_bits_fp),
    .io_deq_bits_branch(fifo_0_io_deq_bits_branch),
    .io_deq_bits_simt_stack(fifo_0_io_deq_bits_simt_stack),
    .io_deq_bits_simt_stack_op(fifo_0_io_deq_bits_simt_stack_op),
    .io_deq_bits_barrier(fifo_0_io_deq_bits_barrier),
    .io_deq_bits_csr(fifo_0_io_deq_bits_csr),
    .io_deq_bits_reverse(fifo_0_io_deq_bits_reverse),
    .io_deq_bits_sel_alu2(fifo_0_io_deq_bits_sel_alu2),
    .io_deq_bits_sel_alu1(fifo_0_io_deq_bits_sel_alu1),
    .io_deq_bits_isvec(fifo_0_io_deq_bits_isvec),
    .io_deq_bits_sel_alu3(fifo_0_io_deq_bits_sel_alu3),
    .io_deq_bits_mask(fifo_0_io_deq_bits_mask),
    .io_deq_bits_sel_imm(fifo_0_io_deq_bits_sel_imm),
    .io_deq_bits_mem_unsigned(fifo_0_io_deq_bits_mem_unsigned),
    .io_deq_bits_alu_fn(fifo_0_io_deq_bits_alu_fn),
    .io_deq_bits_mem(fifo_0_io_deq_bits_mem),
    .io_deq_bits_mem_cmd(fifo_0_io_deq_bits_mem_cmd),
    .io_deq_bits_mop(fifo_0_io_deq_bits_mop),
    .io_deq_bits_reg_idx1(fifo_0_io_deq_bits_reg_idx1),
    .io_deq_bits_reg_idx2(fifo_0_io_deq_bits_reg_idx2),
    .io_deq_bits_reg_idx3(fifo_0_io_deq_bits_reg_idx3),
    .io_deq_bits_reg_idxw(fifo_0_io_deq_bits_reg_idxw),
    .io_deq_bits_wfd(fifo_0_io_deq_bits_wfd),
    .io_deq_bits_fence(fifo_0_io_deq_bits_fence),
    .io_deq_bits_sfu(fifo_0_io_deq_bits_sfu),
    .io_deq_bits_readmask(fifo_0_io_deq_bits_readmask),
    .io_deq_bits_writemask(fifo_0_io_deq_bits_writemask),
    .io_deq_bits_wxd(fifo_0_io_deq_bits_wxd),
    .io_deq_bits_pc(fifo_0_io_deq_bits_pc),
    .io_flush(fifo_0_io_flush)
  );
  QueueWithFlush fifo_1 ( // @[ibuffer.scala 20:24]
    .clock(fifo_1_clock),
    .reset(fifo_1_reset),
    .io_enq_ready(fifo_1_io_enq_ready),
    .io_enq_valid(fifo_1_io_enq_valid),
    .io_enq_bits_inst(fifo_1_io_enq_bits_inst),
    .io_enq_bits_wid(fifo_1_io_enq_bits_wid),
    .io_enq_bits_fp(fifo_1_io_enq_bits_fp),
    .io_enq_bits_branch(fifo_1_io_enq_bits_branch),
    .io_enq_bits_simt_stack(fifo_1_io_enq_bits_simt_stack),
    .io_enq_bits_simt_stack_op(fifo_1_io_enq_bits_simt_stack_op),
    .io_enq_bits_barrier(fifo_1_io_enq_bits_barrier),
    .io_enq_bits_csr(fifo_1_io_enq_bits_csr),
    .io_enq_bits_reverse(fifo_1_io_enq_bits_reverse),
    .io_enq_bits_sel_alu2(fifo_1_io_enq_bits_sel_alu2),
    .io_enq_bits_sel_alu1(fifo_1_io_enq_bits_sel_alu1),
    .io_enq_bits_isvec(fifo_1_io_enq_bits_isvec),
    .io_enq_bits_sel_alu3(fifo_1_io_enq_bits_sel_alu3),
    .io_enq_bits_mask(fifo_1_io_enq_bits_mask),
    .io_enq_bits_sel_imm(fifo_1_io_enq_bits_sel_imm),
    .io_enq_bits_mem_unsigned(fifo_1_io_enq_bits_mem_unsigned),
    .io_enq_bits_alu_fn(fifo_1_io_enq_bits_alu_fn),
    .io_enq_bits_mem(fifo_1_io_enq_bits_mem),
    .io_enq_bits_mem_cmd(fifo_1_io_enq_bits_mem_cmd),
    .io_enq_bits_mop(fifo_1_io_enq_bits_mop),
    .io_enq_bits_reg_idx1(fifo_1_io_enq_bits_reg_idx1),
    .io_enq_bits_reg_idx2(fifo_1_io_enq_bits_reg_idx2),
    .io_enq_bits_reg_idx3(fifo_1_io_enq_bits_reg_idx3),
    .io_enq_bits_reg_idxw(fifo_1_io_enq_bits_reg_idxw),
    .io_enq_bits_wfd(fifo_1_io_enq_bits_wfd),
    .io_enq_bits_fence(fifo_1_io_enq_bits_fence),
    .io_enq_bits_sfu(fifo_1_io_enq_bits_sfu),
    .io_enq_bits_readmask(fifo_1_io_enq_bits_readmask),
    .io_enq_bits_writemask(fifo_1_io_enq_bits_writemask),
    .io_enq_bits_wxd(fifo_1_io_enq_bits_wxd),
    .io_enq_bits_pc(fifo_1_io_enq_bits_pc),
    .io_deq_ready(fifo_1_io_deq_ready),
    .io_deq_valid(fifo_1_io_deq_valid),
    .io_deq_bits_inst(fifo_1_io_deq_bits_inst),
    .io_deq_bits_wid(fifo_1_io_deq_bits_wid),
    .io_deq_bits_fp(fifo_1_io_deq_bits_fp),
    .io_deq_bits_branch(fifo_1_io_deq_bits_branch),
    .io_deq_bits_simt_stack(fifo_1_io_deq_bits_simt_stack),
    .io_deq_bits_simt_stack_op(fifo_1_io_deq_bits_simt_stack_op),
    .io_deq_bits_barrier(fifo_1_io_deq_bits_barrier),
    .io_deq_bits_csr(fifo_1_io_deq_bits_csr),
    .io_deq_bits_reverse(fifo_1_io_deq_bits_reverse),
    .io_deq_bits_sel_alu2(fifo_1_io_deq_bits_sel_alu2),
    .io_deq_bits_sel_alu1(fifo_1_io_deq_bits_sel_alu1),
    .io_deq_bits_isvec(fifo_1_io_deq_bits_isvec),
    .io_deq_bits_sel_alu3(fifo_1_io_deq_bits_sel_alu3),
    .io_deq_bits_mask(fifo_1_io_deq_bits_mask),
    .io_deq_bits_sel_imm(fifo_1_io_deq_bits_sel_imm),
    .io_deq_bits_mem_unsigned(fifo_1_io_deq_bits_mem_unsigned),
    .io_deq_bits_alu_fn(fifo_1_io_deq_bits_alu_fn),
    .io_deq_bits_mem(fifo_1_io_deq_bits_mem),
    .io_deq_bits_mem_cmd(fifo_1_io_deq_bits_mem_cmd),
    .io_deq_bits_mop(fifo_1_io_deq_bits_mop),
    .io_deq_bits_reg_idx1(fifo_1_io_deq_bits_reg_idx1),
    .io_deq_bits_reg_idx2(fifo_1_io_deq_bits_reg_idx2),
    .io_deq_bits_reg_idx3(fifo_1_io_deq_bits_reg_idx3),
    .io_deq_bits_reg_idxw(fifo_1_io_deq_bits_reg_idxw),
    .io_deq_bits_wfd(fifo_1_io_deq_bits_wfd),
    .io_deq_bits_fence(fifo_1_io_deq_bits_fence),
    .io_deq_bits_sfu(fifo_1_io_deq_bits_sfu),
    .io_deq_bits_readmask(fifo_1_io_deq_bits_readmask),
    .io_deq_bits_writemask(fifo_1_io_deq_bits_writemask),
    .io_deq_bits_wxd(fifo_1_io_deq_bits_wxd),
    .io_deq_bits_pc(fifo_1_io_deq_bits_pc),
    .io_flush(fifo_1_io_flush)
  );
  QueueWithFlush fifo_2 ( // @[ibuffer.scala 20:24]
    .clock(fifo_2_clock),
    .reset(fifo_2_reset),
    .io_enq_ready(fifo_2_io_enq_ready),
    .io_enq_valid(fifo_2_io_enq_valid),
    .io_enq_bits_inst(fifo_2_io_enq_bits_inst),
    .io_enq_bits_wid(fifo_2_io_enq_bits_wid),
    .io_enq_bits_fp(fifo_2_io_enq_bits_fp),
    .io_enq_bits_branch(fifo_2_io_enq_bits_branch),
    .io_enq_bits_simt_stack(fifo_2_io_enq_bits_simt_stack),
    .io_enq_bits_simt_stack_op(fifo_2_io_enq_bits_simt_stack_op),
    .io_enq_bits_barrier(fifo_2_io_enq_bits_barrier),
    .io_enq_bits_csr(fifo_2_io_enq_bits_csr),
    .io_enq_bits_reverse(fifo_2_io_enq_bits_reverse),
    .io_enq_bits_sel_alu2(fifo_2_io_enq_bits_sel_alu2),
    .io_enq_bits_sel_alu1(fifo_2_io_enq_bits_sel_alu1),
    .io_enq_bits_isvec(fifo_2_io_enq_bits_isvec),
    .io_enq_bits_sel_alu3(fifo_2_io_enq_bits_sel_alu3),
    .io_enq_bits_mask(fifo_2_io_enq_bits_mask),
    .io_enq_bits_sel_imm(fifo_2_io_enq_bits_sel_imm),
    .io_enq_bits_mem_unsigned(fifo_2_io_enq_bits_mem_unsigned),
    .io_enq_bits_alu_fn(fifo_2_io_enq_bits_alu_fn),
    .io_enq_bits_mem(fifo_2_io_enq_bits_mem),
    .io_enq_bits_mem_cmd(fifo_2_io_enq_bits_mem_cmd),
    .io_enq_bits_mop(fifo_2_io_enq_bits_mop),
    .io_enq_bits_reg_idx1(fifo_2_io_enq_bits_reg_idx1),
    .io_enq_bits_reg_idx2(fifo_2_io_enq_bits_reg_idx2),
    .io_enq_bits_reg_idx3(fifo_2_io_enq_bits_reg_idx3),
    .io_enq_bits_reg_idxw(fifo_2_io_enq_bits_reg_idxw),
    .io_enq_bits_wfd(fifo_2_io_enq_bits_wfd),
    .io_enq_bits_fence(fifo_2_io_enq_bits_fence),
    .io_enq_bits_sfu(fifo_2_io_enq_bits_sfu),
    .io_enq_bits_readmask(fifo_2_io_enq_bits_readmask),
    .io_enq_bits_writemask(fifo_2_io_enq_bits_writemask),
    .io_enq_bits_wxd(fifo_2_io_enq_bits_wxd),
    .io_enq_bits_pc(fifo_2_io_enq_bits_pc),
    .io_deq_ready(fifo_2_io_deq_ready),
    .io_deq_valid(fifo_2_io_deq_valid),
    .io_deq_bits_inst(fifo_2_io_deq_bits_inst),
    .io_deq_bits_wid(fifo_2_io_deq_bits_wid),
    .io_deq_bits_fp(fifo_2_io_deq_bits_fp),
    .io_deq_bits_branch(fifo_2_io_deq_bits_branch),
    .io_deq_bits_simt_stack(fifo_2_io_deq_bits_simt_stack),
    .io_deq_bits_simt_stack_op(fifo_2_io_deq_bits_simt_stack_op),
    .io_deq_bits_barrier(fifo_2_io_deq_bits_barrier),
    .io_deq_bits_csr(fifo_2_io_deq_bits_csr),
    .io_deq_bits_reverse(fifo_2_io_deq_bits_reverse),
    .io_deq_bits_sel_alu2(fifo_2_io_deq_bits_sel_alu2),
    .io_deq_bits_sel_alu1(fifo_2_io_deq_bits_sel_alu1),
    .io_deq_bits_isvec(fifo_2_io_deq_bits_isvec),
    .io_deq_bits_sel_alu3(fifo_2_io_deq_bits_sel_alu3),
    .io_deq_bits_mask(fifo_2_io_deq_bits_mask),
    .io_deq_bits_sel_imm(fifo_2_io_deq_bits_sel_imm),
    .io_deq_bits_mem_unsigned(fifo_2_io_deq_bits_mem_unsigned),
    .io_deq_bits_alu_fn(fifo_2_io_deq_bits_alu_fn),
    .io_deq_bits_mem(fifo_2_io_deq_bits_mem),
    .io_deq_bits_mem_cmd(fifo_2_io_deq_bits_mem_cmd),
    .io_deq_bits_mop(fifo_2_io_deq_bits_mop),
    .io_deq_bits_reg_idx1(fifo_2_io_deq_bits_reg_idx1),
    .io_deq_bits_reg_idx2(fifo_2_io_deq_bits_reg_idx2),
    .io_deq_bits_reg_idx3(fifo_2_io_deq_bits_reg_idx3),
    .io_deq_bits_reg_idxw(fifo_2_io_deq_bits_reg_idxw),
    .io_deq_bits_wfd(fifo_2_io_deq_bits_wfd),
    .io_deq_bits_fence(fifo_2_io_deq_bits_fence),
    .io_deq_bits_sfu(fifo_2_io_deq_bits_sfu),
    .io_deq_bits_readmask(fifo_2_io_deq_bits_readmask),
    .io_deq_bits_writemask(fifo_2_io_deq_bits_writemask),
    .io_deq_bits_wxd(fifo_2_io_deq_bits_wxd),
    .io_deq_bits_pc(fifo_2_io_deq_bits_pc),
    .io_flush(fifo_2_io_flush)
  );
  QueueWithFlush fifo_3 ( // @[ibuffer.scala 20:24]
    .clock(fifo_3_clock),
    .reset(fifo_3_reset),
    .io_enq_ready(fifo_3_io_enq_ready),
    .io_enq_valid(fifo_3_io_enq_valid),
    .io_enq_bits_inst(fifo_3_io_enq_bits_inst),
    .io_enq_bits_wid(fifo_3_io_enq_bits_wid),
    .io_enq_bits_fp(fifo_3_io_enq_bits_fp),
    .io_enq_bits_branch(fifo_3_io_enq_bits_branch),
    .io_enq_bits_simt_stack(fifo_3_io_enq_bits_simt_stack),
    .io_enq_bits_simt_stack_op(fifo_3_io_enq_bits_simt_stack_op),
    .io_enq_bits_barrier(fifo_3_io_enq_bits_barrier),
    .io_enq_bits_csr(fifo_3_io_enq_bits_csr),
    .io_enq_bits_reverse(fifo_3_io_enq_bits_reverse),
    .io_enq_bits_sel_alu2(fifo_3_io_enq_bits_sel_alu2),
    .io_enq_bits_sel_alu1(fifo_3_io_enq_bits_sel_alu1),
    .io_enq_bits_isvec(fifo_3_io_enq_bits_isvec),
    .io_enq_bits_sel_alu3(fifo_3_io_enq_bits_sel_alu3),
    .io_enq_bits_mask(fifo_3_io_enq_bits_mask),
    .io_enq_bits_sel_imm(fifo_3_io_enq_bits_sel_imm),
    .io_enq_bits_mem_unsigned(fifo_3_io_enq_bits_mem_unsigned),
    .io_enq_bits_alu_fn(fifo_3_io_enq_bits_alu_fn),
    .io_enq_bits_mem(fifo_3_io_enq_bits_mem),
    .io_enq_bits_mem_cmd(fifo_3_io_enq_bits_mem_cmd),
    .io_enq_bits_mop(fifo_3_io_enq_bits_mop),
    .io_enq_bits_reg_idx1(fifo_3_io_enq_bits_reg_idx1),
    .io_enq_bits_reg_idx2(fifo_3_io_enq_bits_reg_idx2),
    .io_enq_bits_reg_idx3(fifo_3_io_enq_bits_reg_idx3),
    .io_enq_bits_reg_idxw(fifo_3_io_enq_bits_reg_idxw),
    .io_enq_bits_wfd(fifo_3_io_enq_bits_wfd),
    .io_enq_bits_fence(fifo_3_io_enq_bits_fence),
    .io_enq_bits_sfu(fifo_3_io_enq_bits_sfu),
    .io_enq_bits_readmask(fifo_3_io_enq_bits_readmask),
    .io_enq_bits_writemask(fifo_3_io_enq_bits_writemask),
    .io_enq_bits_wxd(fifo_3_io_enq_bits_wxd),
    .io_enq_bits_pc(fifo_3_io_enq_bits_pc),
    .io_deq_ready(fifo_3_io_deq_ready),
    .io_deq_valid(fifo_3_io_deq_valid),
    .io_deq_bits_inst(fifo_3_io_deq_bits_inst),
    .io_deq_bits_wid(fifo_3_io_deq_bits_wid),
    .io_deq_bits_fp(fifo_3_io_deq_bits_fp),
    .io_deq_bits_branch(fifo_3_io_deq_bits_branch),
    .io_deq_bits_simt_stack(fifo_3_io_deq_bits_simt_stack),
    .io_deq_bits_simt_stack_op(fifo_3_io_deq_bits_simt_stack_op),
    .io_deq_bits_barrier(fifo_3_io_deq_bits_barrier),
    .io_deq_bits_csr(fifo_3_io_deq_bits_csr),
    .io_deq_bits_reverse(fifo_3_io_deq_bits_reverse),
    .io_deq_bits_sel_alu2(fifo_3_io_deq_bits_sel_alu2),
    .io_deq_bits_sel_alu1(fifo_3_io_deq_bits_sel_alu1),
    .io_deq_bits_isvec(fifo_3_io_deq_bits_isvec),
    .io_deq_bits_sel_alu3(fifo_3_io_deq_bits_sel_alu3),
    .io_deq_bits_mask(fifo_3_io_deq_bits_mask),
    .io_deq_bits_sel_imm(fifo_3_io_deq_bits_sel_imm),
    .io_deq_bits_mem_unsigned(fifo_3_io_deq_bits_mem_unsigned),
    .io_deq_bits_alu_fn(fifo_3_io_deq_bits_alu_fn),
    .io_deq_bits_mem(fifo_3_io_deq_bits_mem),
    .io_deq_bits_mem_cmd(fifo_3_io_deq_bits_mem_cmd),
    .io_deq_bits_mop(fifo_3_io_deq_bits_mop),
    .io_deq_bits_reg_idx1(fifo_3_io_deq_bits_reg_idx1),
    .io_deq_bits_reg_idx2(fifo_3_io_deq_bits_reg_idx2),
    .io_deq_bits_reg_idx3(fifo_3_io_deq_bits_reg_idx3),
    .io_deq_bits_reg_idxw(fifo_3_io_deq_bits_reg_idxw),
    .io_deq_bits_wfd(fifo_3_io_deq_bits_wfd),
    .io_deq_bits_fence(fifo_3_io_deq_bits_fence),
    .io_deq_bits_sfu(fifo_3_io_deq_bits_sfu),
    .io_deq_bits_readmask(fifo_3_io_deq_bits_readmask),
    .io_deq_bits_writemask(fifo_3_io_deq_bits_writemask),
    .io_deq_bits_wxd(fifo_3_io_deq_bits_wxd),
    .io_deq_bits_pc(fifo_3_io_deq_bits_pc),
    .io_flush(fifo_3_io_flush)
  );
  assign io_in_ready = _x_single_io_enq_valid_T_6 ? fifo_3_io_enq_ready : _GEN_2; // @[ibuffer.scala 24:{40,52}]
  assign io_out_0_valid = fifo_0_io_deq_valid; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_inst = fifo_0_io_deq_bits_inst; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_wid = fifo_0_io_deq_bits_wid; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_fp = fifo_0_io_deq_bits_fp; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_branch = fifo_0_io_deq_bits_branch; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_simt_stack = fifo_0_io_deq_bits_simt_stack; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_simt_stack_op = fifo_0_io_deq_bits_simt_stack_op; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_barrier = fifo_0_io_deq_bits_barrier; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_csr = fifo_0_io_deq_bits_csr; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_reverse = fifo_0_io_deq_bits_reverse; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_sel_alu2 = fifo_0_io_deq_bits_sel_alu2; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_sel_alu1 = fifo_0_io_deq_bits_sel_alu1; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_isvec = fifo_0_io_deq_bits_isvec; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_sel_alu3 = fifo_0_io_deq_bits_sel_alu3; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_mask = fifo_0_io_deq_bits_mask; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_sel_imm = fifo_0_io_deq_bits_sel_imm; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_mem_unsigned = fifo_0_io_deq_bits_mem_unsigned; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_alu_fn = fifo_0_io_deq_bits_alu_fn; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_mem = fifo_0_io_deq_bits_mem; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_mem_cmd = fifo_0_io_deq_bits_mem_cmd; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_mop = fifo_0_io_deq_bits_mop; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_reg_idx1 = fifo_0_io_deq_bits_reg_idx1; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_reg_idx2 = fifo_0_io_deq_bits_reg_idx2; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_reg_idx3 = fifo_0_io_deq_bits_reg_idx3; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_reg_idxw = fifo_0_io_deq_bits_reg_idxw; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_wfd = fifo_0_io_deq_bits_wfd; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_fence = fifo_0_io_deq_bits_fence; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_sfu = fifo_0_io_deq_bits_sfu; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_readmask = fifo_0_io_deq_bits_readmask; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_writemask = fifo_0_io_deq_bits_writemask; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_wxd = fifo_0_io_deq_bits_wxd; // @[ibuffer.scala 25:16]
  assign io_out_0_bits_pc = fifo_0_io_deq_bits_pc; // @[ibuffer.scala 25:16]
  assign io_out_1_valid = fifo_1_io_deq_valid; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_inst = fifo_1_io_deq_bits_inst; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_wid = fifo_1_io_deq_bits_wid; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_fp = fifo_1_io_deq_bits_fp; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_branch = fifo_1_io_deq_bits_branch; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_simt_stack = fifo_1_io_deq_bits_simt_stack; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_simt_stack_op = fifo_1_io_deq_bits_simt_stack_op; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_barrier = fifo_1_io_deq_bits_barrier; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_csr = fifo_1_io_deq_bits_csr; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_reverse = fifo_1_io_deq_bits_reverse; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_sel_alu2 = fifo_1_io_deq_bits_sel_alu2; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_sel_alu1 = fifo_1_io_deq_bits_sel_alu1; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_isvec = fifo_1_io_deq_bits_isvec; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_sel_alu3 = fifo_1_io_deq_bits_sel_alu3; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_mask = fifo_1_io_deq_bits_mask; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_sel_imm = fifo_1_io_deq_bits_sel_imm; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_mem_unsigned = fifo_1_io_deq_bits_mem_unsigned; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_alu_fn = fifo_1_io_deq_bits_alu_fn; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_mem = fifo_1_io_deq_bits_mem; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_mem_cmd = fifo_1_io_deq_bits_mem_cmd; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_mop = fifo_1_io_deq_bits_mop; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_reg_idx1 = fifo_1_io_deq_bits_reg_idx1; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_reg_idx2 = fifo_1_io_deq_bits_reg_idx2; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_reg_idx3 = fifo_1_io_deq_bits_reg_idx3; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_reg_idxw = fifo_1_io_deq_bits_reg_idxw; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_wfd = fifo_1_io_deq_bits_wfd; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_fence = fifo_1_io_deq_bits_fence; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_sfu = fifo_1_io_deq_bits_sfu; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_readmask = fifo_1_io_deq_bits_readmask; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_writemask = fifo_1_io_deq_bits_writemask; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_wxd = fifo_1_io_deq_bits_wxd; // @[ibuffer.scala 25:16]
  assign io_out_1_bits_pc = fifo_1_io_deq_bits_pc; // @[ibuffer.scala 25:16]
  assign io_out_2_valid = fifo_2_io_deq_valid; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_inst = fifo_2_io_deq_bits_inst; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_wid = fifo_2_io_deq_bits_wid; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_fp = fifo_2_io_deq_bits_fp; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_branch = fifo_2_io_deq_bits_branch; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_simt_stack = fifo_2_io_deq_bits_simt_stack; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_simt_stack_op = fifo_2_io_deq_bits_simt_stack_op; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_barrier = fifo_2_io_deq_bits_barrier; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_csr = fifo_2_io_deq_bits_csr; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_reverse = fifo_2_io_deq_bits_reverse; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_sel_alu2 = fifo_2_io_deq_bits_sel_alu2; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_sel_alu1 = fifo_2_io_deq_bits_sel_alu1; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_isvec = fifo_2_io_deq_bits_isvec; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_sel_alu3 = fifo_2_io_deq_bits_sel_alu3; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_mask = fifo_2_io_deq_bits_mask; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_sel_imm = fifo_2_io_deq_bits_sel_imm; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_mem_unsigned = fifo_2_io_deq_bits_mem_unsigned; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_alu_fn = fifo_2_io_deq_bits_alu_fn; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_mem = fifo_2_io_deq_bits_mem; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_mem_cmd = fifo_2_io_deq_bits_mem_cmd; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_mop = fifo_2_io_deq_bits_mop; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_reg_idx1 = fifo_2_io_deq_bits_reg_idx1; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_reg_idx2 = fifo_2_io_deq_bits_reg_idx2; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_reg_idx3 = fifo_2_io_deq_bits_reg_idx3; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_reg_idxw = fifo_2_io_deq_bits_reg_idxw; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_wfd = fifo_2_io_deq_bits_wfd; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_fence = fifo_2_io_deq_bits_fence; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_sfu = fifo_2_io_deq_bits_sfu; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_readmask = fifo_2_io_deq_bits_readmask; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_writemask = fifo_2_io_deq_bits_writemask; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_wxd = fifo_2_io_deq_bits_wxd; // @[ibuffer.scala 25:16]
  assign io_out_2_bits_pc = fifo_2_io_deq_bits_pc; // @[ibuffer.scala 25:16]
  assign io_out_3_valid = fifo_3_io_deq_valid; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_inst = fifo_3_io_deq_bits_inst; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_wid = fifo_3_io_deq_bits_wid; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_fp = fifo_3_io_deq_bits_fp; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_branch = fifo_3_io_deq_bits_branch; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_simt_stack = fifo_3_io_deq_bits_simt_stack; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_simt_stack_op = fifo_3_io_deq_bits_simt_stack_op; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_barrier = fifo_3_io_deq_bits_barrier; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_csr = fifo_3_io_deq_bits_csr; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_reverse = fifo_3_io_deq_bits_reverse; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_sel_alu2 = fifo_3_io_deq_bits_sel_alu2; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_sel_alu1 = fifo_3_io_deq_bits_sel_alu1; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_isvec = fifo_3_io_deq_bits_isvec; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_sel_alu3 = fifo_3_io_deq_bits_sel_alu3; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_mask = fifo_3_io_deq_bits_mask; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_sel_imm = fifo_3_io_deq_bits_sel_imm; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_mem_unsigned = fifo_3_io_deq_bits_mem_unsigned; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_alu_fn = fifo_3_io_deq_bits_alu_fn; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_mem = fifo_3_io_deq_bits_mem; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_mem_cmd = fifo_3_io_deq_bits_mem_cmd; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_mop = fifo_3_io_deq_bits_mop; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_reg_idx1 = fifo_3_io_deq_bits_reg_idx1; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_reg_idx2 = fifo_3_io_deq_bits_reg_idx2; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_reg_idx3 = fifo_3_io_deq_bits_reg_idx3; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_reg_idxw = fifo_3_io_deq_bits_reg_idxw; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_wfd = fifo_3_io_deq_bits_wfd; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_fence = fifo_3_io_deq_bits_fence; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_sfu = fifo_3_io_deq_bits_sfu; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_readmask = fifo_3_io_deq_bits_readmask; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_writemask = fifo_3_io_deq_bits_writemask; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_wxd = fifo_3_io_deq_bits_wxd; // @[ibuffer.scala 25:16]
  assign io_out_3_bits_pc = fifo_3_io_deq_bits_pc; // @[ibuffer.scala 25:16]
  assign io_ibuffer_ready_0 = fifo_0_io_enq_ready; // @[ibuffer.scala 21:26]
  assign io_ibuffer_ready_1 = fifo_1_io_enq_ready; // @[ibuffer.scala 21:26]
  assign io_ibuffer_ready_2 = fifo_2_io_enq_ready; // @[ibuffer.scala 21:26]
  assign io_ibuffer_ready_3 = fifo_3_io_enq_ready; // @[ibuffer.scala 21:26]
  assign fifo_0_clock = clock;
  assign fifo_0_reset = reset;
  assign fifo_0_io_enq_valid = 2'h0 == io_in_bits_wid & io_in_valid; // @[ibuffer.scala 23:33]
  assign fifo_0_io_enq_bits_inst = io_in_bits_inst; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_wid = io_in_bits_wid; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_fp = io_in_bits_fp; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_branch = io_in_bits_branch; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_simt_stack = io_in_bits_simt_stack; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_simt_stack_op = io_in_bits_simt_stack_op; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_barrier = io_in_bits_barrier; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_csr = io_in_bits_csr; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_reverse = io_in_bits_reverse; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_sel_alu2 = io_in_bits_sel_alu2; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_sel_alu1 = io_in_bits_sel_alu1; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_isvec = io_in_bits_isvec; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_sel_alu3 = io_in_bits_sel_alu3; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_mask = io_in_bits_mask; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_sel_imm = io_in_bits_sel_imm; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_mem_unsigned = io_in_bits_mem_unsigned; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_alu_fn = io_in_bits_alu_fn; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_mem = io_in_bits_mem; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_mem_cmd = io_in_bits_mem_cmd; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_mop = io_in_bits_mop; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_reg_idx1 = io_in_bits_reg_idx1; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_reg_idx2 = io_in_bits_reg_idx2; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_reg_idx3 = io_in_bits_reg_idx3; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_reg_idxw = io_in_bits_reg_idxw; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_wfd = io_in_bits_wfd; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_fence = io_in_bits_fence; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_sfu = io_in_bits_sfu; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_readmask = io_in_bits_readmask; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_writemask = io_in_bits_writemask; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_wxd = io_in_bits_wxd; // @[ibuffer.scala 22:27]
  assign fifo_0_io_enq_bits_pc = io_in_bits_pc; // @[ibuffer.scala 22:27]
  assign fifo_0_io_deq_ready = io_out_0_ready; // @[ibuffer.scala 25:16]
  assign fifo_0_io_flush = io_flush_valid & 2'h0 == io_flush_bits; // @[ibuffer.scala 26:37]
  assign fifo_1_clock = clock;
  assign fifo_1_reset = reset;
  assign fifo_1_io_enq_valid = 2'h1 == io_in_bits_wid & io_in_valid; // @[ibuffer.scala 23:33]
  assign fifo_1_io_enq_bits_inst = io_in_bits_inst; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_wid = io_in_bits_wid; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_fp = io_in_bits_fp; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_branch = io_in_bits_branch; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_simt_stack = io_in_bits_simt_stack; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_simt_stack_op = io_in_bits_simt_stack_op; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_barrier = io_in_bits_barrier; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_csr = io_in_bits_csr; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_reverse = io_in_bits_reverse; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_sel_alu2 = io_in_bits_sel_alu2; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_sel_alu1 = io_in_bits_sel_alu1; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_isvec = io_in_bits_isvec; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_sel_alu3 = io_in_bits_sel_alu3; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_mask = io_in_bits_mask; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_sel_imm = io_in_bits_sel_imm; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_mem_unsigned = io_in_bits_mem_unsigned; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_alu_fn = io_in_bits_alu_fn; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_mem = io_in_bits_mem; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_mem_cmd = io_in_bits_mem_cmd; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_mop = io_in_bits_mop; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_reg_idx1 = io_in_bits_reg_idx1; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_reg_idx2 = io_in_bits_reg_idx2; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_reg_idx3 = io_in_bits_reg_idx3; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_reg_idxw = io_in_bits_reg_idxw; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_wfd = io_in_bits_wfd; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_fence = io_in_bits_fence; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_sfu = io_in_bits_sfu; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_readmask = io_in_bits_readmask; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_writemask = io_in_bits_writemask; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_wxd = io_in_bits_wxd; // @[ibuffer.scala 22:27]
  assign fifo_1_io_enq_bits_pc = io_in_bits_pc; // @[ibuffer.scala 22:27]
  assign fifo_1_io_deq_ready = io_out_1_ready; // @[ibuffer.scala 25:16]
  assign fifo_1_io_flush = io_flush_valid & 2'h1 == io_flush_bits; // @[ibuffer.scala 26:37]
  assign fifo_2_clock = clock;
  assign fifo_2_reset = reset;
  assign fifo_2_io_enq_valid = 2'h2 == io_in_bits_wid & io_in_valid; // @[ibuffer.scala 23:33]
  assign fifo_2_io_enq_bits_inst = io_in_bits_inst; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_wid = io_in_bits_wid; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_fp = io_in_bits_fp; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_branch = io_in_bits_branch; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_simt_stack = io_in_bits_simt_stack; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_simt_stack_op = io_in_bits_simt_stack_op; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_barrier = io_in_bits_barrier; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_csr = io_in_bits_csr; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_reverse = io_in_bits_reverse; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_sel_alu2 = io_in_bits_sel_alu2; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_sel_alu1 = io_in_bits_sel_alu1; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_isvec = io_in_bits_isvec; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_sel_alu3 = io_in_bits_sel_alu3; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_mask = io_in_bits_mask; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_sel_imm = io_in_bits_sel_imm; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_mem_unsigned = io_in_bits_mem_unsigned; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_alu_fn = io_in_bits_alu_fn; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_mem = io_in_bits_mem; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_mem_cmd = io_in_bits_mem_cmd; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_mop = io_in_bits_mop; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_reg_idx1 = io_in_bits_reg_idx1; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_reg_idx2 = io_in_bits_reg_idx2; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_reg_idx3 = io_in_bits_reg_idx3; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_reg_idxw = io_in_bits_reg_idxw; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_wfd = io_in_bits_wfd; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_fence = io_in_bits_fence; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_sfu = io_in_bits_sfu; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_readmask = io_in_bits_readmask; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_writemask = io_in_bits_writemask; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_wxd = io_in_bits_wxd; // @[ibuffer.scala 22:27]
  assign fifo_2_io_enq_bits_pc = io_in_bits_pc; // @[ibuffer.scala 22:27]
  assign fifo_2_io_deq_ready = io_out_2_ready; // @[ibuffer.scala 25:16]
  assign fifo_2_io_flush = io_flush_valid & 2'h2 == io_flush_bits; // @[ibuffer.scala 26:37]
  assign fifo_3_clock = clock;
  assign fifo_3_reset = reset;
  assign fifo_3_io_enq_valid = 2'h3 == io_in_bits_wid & io_in_valid; // @[ibuffer.scala 23:33]
  assign fifo_3_io_enq_bits_inst = io_in_bits_inst; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_wid = io_in_bits_wid; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_fp = io_in_bits_fp; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_branch = io_in_bits_branch; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_simt_stack = io_in_bits_simt_stack; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_simt_stack_op = io_in_bits_simt_stack_op; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_barrier = io_in_bits_barrier; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_csr = io_in_bits_csr; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_reverse = io_in_bits_reverse; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_sel_alu2 = io_in_bits_sel_alu2; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_sel_alu1 = io_in_bits_sel_alu1; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_isvec = io_in_bits_isvec; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_sel_alu3 = io_in_bits_sel_alu3; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_mask = io_in_bits_mask; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_sel_imm = io_in_bits_sel_imm; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_mem_unsigned = io_in_bits_mem_unsigned; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_alu_fn = io_in_bits_alu_fn; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_mem = io_in_bits_mem; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_mem_cmd = io_in_bits_mem_cmd; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_mop = io_in_bits_mop; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_reg_idx1 = io_in_bits_reg_idx1; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_reg_idx2 = io_in_bits_reg_idx2; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_reg_idx3 = io_in_bits_reg_idx3; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_reg_idxw = io_in_bits_reg_idxw; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_wfd = io_in_bits_wfd; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_fence = io_in_bits_fence; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_sfu = io_in_bits_sfu; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_readmask = io_in_bits_readmask; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_writemask = io_in_bits_writemask; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_wxd = io_in_bits_wxd; // @[ibuffer.scala 22:27]
  assign fifo_3_io_enq_bits_pc = io_in_bits_pc; // @[ibuffer.scala 22:27]
  assign fifo_3_io_deq_ready = io_out_3_ready; // @[ibuffer.scala 25:16]
  assign fifo_3_io_flush = io_flush_valid & 2'h3 == io_flush_bits; // @[ibuffer.scala 26:37]
endmodule
module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_inst,
  input  [1:0]  io_in_0_bits_wid,
  input         io_in_0_bits_fp,
  input  [1:0]  io_in_0_bits_branch,
  input         io_in_0_bits_simt_stack,
  input         io_in_0_bits_simt_stack_op,
  input         io_in_0_bits_barrier,
  input  [1:0]  io_in_0_bits_csr,
  input         io_in_0_bits_reverse,
  input  [1:0]  io_in_0_bits_sel_alu2,
  input  [1:0]  io_in_0_bits_sel_alu1,
  input         io_in_0_bits_isvec,
  input  [1:0]  io_in_0_bits_sel_alu3,
  input         io_in_0_bits_mask,
  input  [2:0]  io_in_0_bits_sel_imm,
  input         io_in_0_bits_mem_unsigned,
  input  [5:0]  io_in_0_bits_alu_fn,
  input         io_in_0_bits_mem,
  input  [1:0]  io_in_0_bits_mem_cmd,
  input  [1:0]  io_in_0_bits_mop,
  input  [4:0]  io_in_0_bits_reg_idx1,
  input  [4:0]  io_in_0_bits_reg_idx2,
  input  [4:0]  io_in_0_bits_reg_idx3,
  input  [4:0]  io_in_0_bits_reg_idxw,
  input         io_in_0_bits_wfd,
  input         io_in_0_bits_fence,
  input         io_in_0_bits_sfu,
  input         io_in_0_bits_readmask,
  input         io_in_0_bits_writemask,
  input         io_in_0_bits_wxd,
  input  [31:0] io_in_0_bits_pc,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_inst,
  input  [1:0]  io_in_1_bits_wid,
  input         io_in_1_bits_fp,
  input  [1:0]  io_in_1_bits_branch,
  input         io_in_1_bits_simt_stack,
  input         io_in_1_bits_simt_stack_op,
  input         io_in_1_bits_barrier,
  input  [1:0]  io_in_1_bits_csr,
  input         io_in_1_bits_reverse,
  input  [1:0]  io_in_1_bits_sel_alu2,
  input  [1:0]  io_in_1_bits_sel_alu1,
  input         io_in_1_bits_isvec,
  input  [1:0]  io_in_1_bits_sel_alu3,
  input         io_in_1_bits_mask,
  input  [2:0]  io_in_1_bits_sel_imm,
  input         io_in_1_bits_mem_unsigned,
  input  [5:0]  io_in_1_bits_alu_fn,
  input         io_in_1_bits_mem,
  input  [1:0]  io_in_1_bits_mem_cmd,
  input  [1:0]  io_in_1_bits_mop,
  input  [4:0]  io_in_1_bits_reg_idx1,
  input  [4:0]  io_in_1_bits_reg_idx2,
  input  [4:0]  io_in_1_bits_reg_idx3,
  input  [4:0]  io_in_1_bits_reg_idxw,
  input         io_in_1_bits_wfd,
  input         io_in_1_bits_fence,
  input         io_in_1_bits_sfu,
  input         io_in_1_bits_readmask,
  input         io_in_1_bits_writemask,
  input         io_in_1_bits_wxd,
  input  [31:0] io_in_1_bits_pc,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_inst,
  input  [1:0]  io_in_2_bits_wid,
  input         io_in_2_bits_fp,
  input  [1:0]  io_in_2_bits_branch,
  input         io_in_2_bits_simt_stack,
  input         io_in_2_bits_simt_stack_op,
  input         io_in_2_bits_barrier,
  input  [1:0]  io_in_2_bits_csr,
  input         io_in_2_bits_reverse,
  input  [1:0]  io_in_2_bits_sel_alu2,
  input  [1:0]  io_in_2_bits_sel_alu1,
  input         io_in_2_bits_isvec,
  input  [1:0]  io_in_2_bits_sel_alu3,
  input         io_in_2_bits_mask,
  input  [2:0]  io_in_2_bits_sel_imm,
  input         io_in_2_bits_mem_unsigned,
  input  [5:0]  io_in_2_bits_alu_fn,
  input         io_in_2_bits_mem,
  input  [1:0]  io_in_2_bits_mem_cmd,
  input  [1:0]  io_in_2_bits_mop,
  input  [4:0]  io_in_2_bits_reg_idx1,
  input  [4:0]  io_in_2_bits_reg_idx2,
  input  [4:0]  io_in_2_bits_reg_idx3,
  input  [4:0]  io_in_2_bits_reg_idxw,
  input         io_in_2_bits_wfd,
  input         io_in_2_bits_fence,
  input         io_in_2_bits_sfu,
  input         io_in_2_bits_readmask,
  input         io_in_2_bits_writemask,
  input         io_in_2_bits_wxd,
  input  [31:0] io_in_2_bits_pc,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_inst,
  input  [1:0]  io_in_3_bits_wid,
  input         io_in_3_bits_fp,
  input  [1:0]  io_in_3_bits_branch,
  input         io_in_3_bits_simt_stack,
  input         io_in_3_bits_simt_stack_op,
  input         io_in_3_bits_barrier,
  input  [1:0]  io_in_3_bits_csr,
  input         io_in_3_bits_reverse,
  input  [1:0]  io_in_3_bits_sel_alu2,
  input  [1:0]  io_in_3_bits_sel_alu1,
  input         io_in_3_bits_isvec,
  input  [1:0]  io_in_3_bits_sel_alu3,
  input         io_in_3_bits_mask,
  input  [2:0]  io_in_3_bits_sel_imm,
  input         io_in_3_bits_mem_unsigned,
  input  [5:0]  io_in_3_bits_alu_fn,
  input         io_in_3_bits_mem,
  input  [1:0]  io_in_3_bits_mem_cmd,
  input  [1:0]  io_in_3_bits_mop,
  input  [4:0]  io_in_3_bits_reg_idx1,
  input  [4:0]  io_in_3_bits_reg_idx2,
  input  [4:0]  io_in_3_bits_reg_idx3,
  input  [4:0]  io_in_3_bits_reg_idxw,
  input         io_in_3_bits_wfd,
  input         io_in_3_bits_fence,
  input         io_in_3_bits_sfu,
  input         io_in_3_bits_readmask,
  input         io_in_3_bits_writemask,
  input         io_in_3_bits_wxd,
  input  [31:0] io_in_3_bits_pc,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_inst,
  output [1:0]  io_out_bits_wid,
  output        io_out_bits_fp,
  output [1:0]  io_out_bits_branch,
  output        io_out_bits_simt_stack,
  output        io_out_bits_simt_stack_op,
  output        io_out_bits_barrier,
  output [1:0]  io_out_bits_csr,
  output        io_out_bits_reverse,
  output [1:0]  io_out_bits_sel_alu2,
  output [1:0]  io_out_bits_sel_alu1,
  output        io_out_bits_isvec,
  output [1:0]  io_out_bits_sel_alu3,
  output        io_out_bits_mask,
  output [2:0]  io_out_bits_sel_imm,
  output        io_out_bits_mem_unsigned,
  output [5:0]  io_out_bits_alu_fn,
  output        io_out_bits_mem,
  output [1:0]  io_out_bits_mem_cmd,
  output [1:0]  io_out_bits_mop,
  output [4:0]  io_out_bits_reg_idx1,
  output [4:0]  io_out_bits_reg_idx2,
  output [4:0]  io_out_bits_reg_idx3,
  output [4:0]  io_out_bits_reg_idxw,
  output        io_out_bits_wfd,
  output        io_out_bits_fence,
  output        io_out_bits_sfu,
  output        io_out_bits_readmask,
  output        io_out_bits_writemask,
  output        io_out_bits_wxd,
  output [31:0] io_out_bits_pc,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 56:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 56:{16,16}]
  wire [31:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_pc : io_in_0_bits_pc; // @[Arbiter.scala 57:{15,15}]
  wire [31:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_pc : _GEN_5; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_wxd : io_in_0_bits_wxd; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_10 = 2'h2 == io_chosen ? io_in_2_bits_wxd : _GEN_9; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_writemask : io_in_0_bits_writemask; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_writemask : _GEN_13; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_readmask : io_in_0_bits_readmask; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_readmask : _GEN_17; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_sfu : io_in_0_bits_sfu; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_sfu : _GEN_21; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_25 = 2'h1 == io_chosen ? io_in_1_bits_fence : io_in_0_bits_fence; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_fence : _GEN_25; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_29 = 2'h1 == io_chosen ? io_in_1_bits_wfd : io_in_0_bits_wfd; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_30 = 2'h2 == io_chosen ? io_in_2_bits_wfd : _GEN_29; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_33 = 2'h1 == io_chosen ? io_in_1_bits_reg_idxw : io_in_0_bits_reg_idxw; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_reg_idxw : _GEN_33; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_37 = 2'h1 == io_chosen ? io_in_1_bits_reg_idx3 : io_in_0_bits_reg_idx3; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_38 = 2'h2 == io_chosen ? io_in_2_bits_reg_idx3 : _GEN_37; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_41 = 2'h1 == io_chosen ? io_in_1_bits_reg_idx2 : io_in_0_bits_reg_idx2; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_42 = 2'h2 == io_chosen ? io_in_2_bits_reg_idx2 : _GEN_41; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_45 = 2'h1 == io_chosen ? io_in_1_bits_reg_idx1 : io_in_0_bits_reg_idx1; // @[Arbiter.scala 57:{15,15}]
  wire [4:0] _GEN_46 = 2'h2 == io_chosen ? io_in_2_bits_reg_idx1 : _GEN_45; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_49 = 2'h1 == io_chosen ? io_in_1_bits_mop : io_in_0_bits_mop; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_50 = 2'h2 == io_chosen ? io_in_2_bits_mop : _GEN_49; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_53 = 2'h1 == io_chosen ? io_in_1_bits_mem_cmd : io_in_0_bits_mem_cmd; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_54 = 2'h2 == io_chosen ? io_in_2_bits_mem_cmd : _GEN_53; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_57 = 2'h1 == io_chosen ? io_in_1_bits_mem : io_in_0_bits_mem; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_58 = 2'h2 == io_chosen ? io_in_2_bits_mem : _GEN_57; // @[Arbiter.scala 57:{15,15}]
  wire [5:0] _GEN_61 = 2'h1 == io_chosen ? io_in_1_bits_alu_fn : io_in_0_bits_alu_fn; // @[Arbiter.scala 57:{15,15}]
  wire [5:0] _GEN_62 = 2'h2 == io_chosen ? io_in_2_bits_alu_fn : _GEN_61; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_65 = 2'h1 == io_chosen ? io_in_1_bits_mem_unsigned : io_in_0_bits_mem_unsigned; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_66 = 2'h2 == io_chosen ? io_in_2_bits_mem_unsigned : _GEN_65; // @[Arbiter.scala 57:{15,15}]
  wire [2:0] _GEN_73 = 2'h1 == io_chosen ? io_in_1_bits_sel_imm : io_in_0_bits_sel_imm; // @[Arbiter.scala 57:{15,15}]
  wire [2:0] _GEN_74 = 2'h2 == io_chosen ? io_in_2_bits_sel_imm : _GEN_73; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_77 = 2'h1 == io_chosen ? io_in_1_bits_mask : io_in_0_bits_mask; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_78 = 2'h2 == io_chosen ? io_in_2_bits_mask : _GEN_77; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_81 = 2'h1 == io_chosen ? io_in_1_bits_sel_alu3 : io_in_0_bits_sel_alu3; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_82 = 2'h2 == io_chosen ? io_in_2_bits_sel_alu3 : _GEN_81; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_85 = 2'h1 == io_chosen ? io_in_1_bits_isvec : io_in_0_bits_isvec; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_86 = 2'h2 == io_chosen ? io_in_2_bits_isvec : _GEN_85; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_89 = 2'h1 == io_chosen ? io_in_1_bits_sel_alu1 : io_in_0_bits_sel_alu1; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_90 = 2'h2 == io_chosen ? io_in_2_bits_sel_alu1 : _GEN_89; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_93 = 2'h1 == io_chosen ? io_in_1_bits_sel_alu2 : io_in_0_bits_sel_alu2; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_94 = 2'h2 == io_chosen ? io_in_2_bits_sel_alu2 : _GEN_93; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_97 = 2'h1 == io_chosen ? io_in_1_bits_reverse : io_in_0_bits_reverse; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_98 = 2'h2 == io_chosen ? io_in_2_bits_reverse : _GEN_97; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_101 = 2'h1 == io_chosen ? io_in_1_bits_csr : io_in_0_bits_csr; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_102 = 2'h2 == io_chosen ? io_in_2_bits_csr : _GEN_101; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_105 = 2'h1 == io_chosen ? io_in_1_bits_barrier : io_in_0_bits_barrier; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_106 = 2'h2 == io_chosen ? io_in_2_bits_barrier : _GEN_105; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_109 = 2'h1 == io_chosen ? io_in_1_bits_simt_stack_op : io_in_0_bits_simt_stack_op; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_110 = 2'h2 == io_chosen ? io_in_2_bits_simt_stack_op : _GEN_109; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_113 = 2'h1 == io_chosen ? io_in_1_bits_simt_stack : io_in_0_bits_simt_stack; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_114 = 2'h2 == io_chosen ? io_in_2_bits_simt_stack : _GEN_113; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_117 = 2'h1 == io_chosen ? io_in_1_bits_branch : io_in_0_bits_branch; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_118 = 2'h2 == io_chosen ? io_in_2_bits_branch : _GEN_117; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_121 = 2'h1 == io_chosen ? io_in_1_bits_fp : io_in_0_bits_fp; // @[Arbiter.scala 57:{15,15}]
  wire  _GEN_122 = 2'h2 == io_chosen ? io_in_2_bits_fp : _GEN_121; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_125 = 2'h1 == io_chosen ? io_in_1_bits_wid : io_in_0_bits_wid; // @[Arbiter.scala 57:{15,15}]
  wire [1:0] _GEN_126 = 2'h2 == io_chosen ? io_in_2_bits_wid : _GEN_125; // @[Arbiter.scala 57:{15,15}]
  wire [31:0] _GEN_129 = 2'h1 == io_chosen ? io_in_1_bits_inst : io_in_0_bits_inst; // @[Arbiter.scala 57:{15,15}]
  wire [31:0] _GEN_130 = 2'h2 == io_chosen ? io_in_2_bits_inst : _GEN_129; // @[Arbiter.scala 57:{15,15}]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 50:35]
  reg [1:0] lastGrant; // @[Reg.scala 16:16]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbiter.scala 82:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbiter.scala 82:49]
  wire  grantMask_3 = 2'h3 > lastGrant; // @[Arbiter.scala 82:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 83:76]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 83:76]
  wire  validMask_3 = io_in_3_valid & grantMask_3; // @[Arbiter.scala 83:76]
  wire  ctrl_2 = ~validMask_1; // @[Arbiter.scala 46:78]
  wire  ctrl_3 = ~(validMask_1 | validMask_2); // @[Arbiter.scala 46:78]
  wire  ctrl_4 = ~(validMask_1 | validMask_2 | validMask_3); // @[Arbiter.scala 46:78]
  wire  ctrl_5 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid); // @[Arbiter.scala 46:78]
  wire  ctrl_6 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 46:78]
  wire  ctrl_7 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 46:78]
  wire  _T_3 = grantMask_1 | ctrl_5; // @[Arbiter.scala 87:50]
  wire  _T_5 = ctrl_2 & grantMask_2 | ctrl_6; // @[Arbiter.scala 87:50]
  wire  _T_7 = ctrl_3 & grantMask_3 | ctrl_7; // @[Arbiter.scala 87:50]
  wire [1:0] _GEN_133 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 92:{26,35}]
  wire [1:0] _GEN_134 = io_in_1_valid ? 2'h1 : _GEN_133; // @[Arbiter.scala 92:{26,35}]
  wire [1:0] _GEN_135 = io_in_0_valid ? 2'h0 : _GEN_134; // @[Arbiter.scala 92:{26,35}]
  wire [1:0] _GEN_136 = validMask_3 ? 2'h3 : _GEN_135; // @[Arbiter.scala 94:{24,33}]
  wire [1:0] _GEN_137 = validMask_2 ? 2'h2 : _GEN_136; // @[Arbiter.scala 94:{24,33}]
  assign io_in_0_ready = ctrl_4 & io_out_ready; // @[Arbiter.scala 75:21]
  assign io_in_1_ready = _T_3 & io_out_ready; // @[Arbiter.scala 75:21]
  assign io_in_2_ready = _T_5 & io_out_ready; // @[Arbiter.scala 75:21]
  assign io_in_3_ready = _T_7 & io_out_ready; // @[Arbiter.scala 75:21]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 56:{16,16}]
  assign io_out_bits_inst = 2'h3 == io_chosen ? io_in_3_bits_inst : _GEN_130; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_wid = 2'h3 == io_chosen ? io_in_3_bits_wid : _GEN_126; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_fp = 2'h3 == io_chosen ? io_in_3_bits_fp : _GEN_122; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_branch = 2'h3 == io_chosen ? io_in_3_bits_branch : _GEN_118; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_simt_stack = 2'h3 == io_chosen ? io_in_3_bits_simt_stack : _GEN_114; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_simt_stack_op = 2'h3 == io_chosen ? io_in_3_bits_simt_stack_op : _GEN_110; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_barrier = 2'h3 == io_chosen ? io_in_3_bits_barrier : _GEN_106; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_csr = 2'h3 == io_chosen ? io_in_3_bits_csr : _GEN_102; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_reverse = 2'h3 == io_chosen ? io_in_3_bits_reverse : _GEN_98; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_sel_alu2 = 2'h3 == io_chosen ? io_in_3_bits_sel_alu2 : _GEN_94; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_sel_alu1 = 2'h3 == io_chosen ? io_in_3_bits_sel_alu1 : _GEN_90; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_isvec = 2'h3 == io_chosen ? io_in_3_bits_isvec : _GEN_86; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_sel_alu3 = 2'h3 == io_chosen ? io_in_3_bits_sel_alu3 : _GEN_82; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_mask = 2'h3 == io_chosen ? io_in_3_bits_mask : _GEN_78; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_sel_imm = 2'h3 == io_chosen ? io_in_3_bits_sel_imm : _GEN_74; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_mem_unsigned = 2'h3 == io_chosen ? io_in_3_bits_mem_unsigned : _GEN_66; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_alu_fn = 2'h3 == io_chosen ? io_in_3_bits_alu_fn : _GEN_62; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_mem = 2'h3 == io_chosen ? io_in_3_bits_mem : _GEN_58; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_mem_cmd = 2'h3 == io_chosen ? io_in_3_bits_mem_cmd : _GEN_54; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_mop = 2'h3 == io_chosen ? io_in_3_bits_mop : _GEN_50; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_reg_idx1 = 2'h3 == io_chosen ? io_in_3_bits_reg_idx1 : _GEN_46; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_reg_idx2 = 2'h3 == io_chosen ? io_in_3_bits_reg_idx2 : _GEN_42; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_reg_idx3 = 2'h3 == io_chosen ? io_in_3_bits_reg_idx3 : _GEN_38; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_reg_idxw = 2'h3 == io_chosen ? io_in_3_bits_reg_idxw : _GEN_34; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_wfd = 2'h3 == io_chosen ? io_in_3_bits_wfd : _GEN_30; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_fence = 2'h3 == io_chosen ? io_in_3_bits_fence : _GEN_26; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_sfu = 2'h3 == io_chosen ? io_in_3_bits_sfu : _GEN_22; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_readmask = 2'h3 == io_chosen ? io_in_3_bits_readmask : _GEN_18; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_writemask = 2'h3 == io_chosen ? io_in_3_bits_writemask : _GEN_14; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_wxd = 2'h3 == io_chosen ? io_in_3_bits_wxd : _GEN_10; // @[Arbiter.scala 57:{15,15}]
  assign io_out_bits_pc = 2'h3 == io_chosen ? io_in_3_bits_pc : _GEN_6; // @[Arbiter.scala 57:{15,15}]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_137; // @[Arbiter.scala 94:{24,33}]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 17:18]
      lastGrant <= io_chosen; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ibuffer2issue(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_inst,
  input  [1:0]  io_in_0_bits_wid,
  input         io_in_0_bits_fp,
  input  [1:0]  io_in_0_bits_branch,
  input         io_in_0_bits_simt_stack,
  input         io_in_0_bits_simt_stack_op,
  input         io_in_0_bits_barrier,
  input  [1:0]  io_in_0_bits_csr,
  input         io_in_0_bits_reverse,
  input  [1:0]  io_in_0_bits_sel_alu2,
  input  [1:0]  io_in_0_bits_sel_alu1,
  input         io_in_0_bits_isvec,
  input  [1:0]  io_in_0_bits_sel_alu3,
  input         io_in_0_bits_mask,
  input  [2:0]  io_in_0_bits_sel_imm,
  input         io_in_0_bits_mem_unsigned,
  input  [5:0]  io_in_0_bits_alu_fn,
  input         io_in_0_bits_mem,
  input  [1:0]  io_in_0_bits_mem_cmd,
  input  [1:0]  io_in_0_bits_mop,
  input  [4:0]  io_in_0_bits_reg_idx1,
  input  [4:0]  io_in_0_bits_reg_idx2,
  input  [4:0]  io_in_0_bits_reg_idx3,
  input  [4:0]  io_in_0_bits_reg_idxw,
  input         io_in_0_bits_wfd,
  input         io_in_0_bits_fence,
  input         io_in_0_bits_sfu,
  input         io_in_0_bits_readmask,
  input         io_in_0_bits_writemask,
  input         io_in_0_bits_wxd,
  input  [31:0] io_in_0_bits_pc,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_inst,
  input  [1:0]  io_in_1_bits_wid,
  input         io_in_1_bits_fp,
  input  [1:0]  io_in_1_bits_branch,
  input         io_in_1_bits_simt_stack,
  input         io_in_1_bits_simt_stack_op,
  input         io_in_1_bits_barrier,
  input  [1:0]  io_in_1_bits_csr,
  input         io_in_1_bits_reverse,
  input  [1:0]  io_in_1_bits_sel_alu2,
  input  [1:0]  io_in_1_bits_sel_alu1,
  input         io_in_1_bits_isvec,
  input  [1:0]  io_in_1_bits_sel_alu3,
  input         io_in_1_bits_mask,
  input  [2:0]  io_in_1_bits_sel_imm,
  input         io_in_1_bits_mem_unsigned,
  input  [5:0]  io_in_1_bits_alu_fn,
  input         io_in_1_bits_mem,
  input  [1:0]  io_in_1_bits_mem_cmd,
  input  [1:0]  io_in_1_bits_mop,
  input  [4:0]  io_in_1_bits_reg_idx1,
  input  [4:0]  io_in_1_bits_reg_idx2,
  input  [4:0]  io_in_1_bits_reg_idx3,
  input  [4:0]  io_in_1_bits_reg_idxw,
  input         io_in_1_bits_wfd,
  input         io_in_1_bits_fence,
  input         io_in_1_bits_sfu,
  input         io_in_1_bits_readmask,
  input         io_in_1_bits_writemask,
  input         io_in_1_bits_wxd,
  input  [31:0] io_in_1_bits_pc,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_inst,
  input  [1:0]  io_in_2_bits_wid,
  input         io_in_2_bits_fp,
  input  [1:0]  io_in_2_bits_branch,
  input         io_in_2_bits_simt_stack,
  input         io_in_2_bits_simt_stack_op,
  input         io_in_2_bits_barrier,
  input  [1:0]  io_in_2_bits_csr,
  input         io_in_2_bits_reverse,
  input  [1:0]  io_in_2_bits_sel_alu2,
  input  [1:0]  io_in_2_bits_sel_alu1,
  input         io_in_2_bits_isvec,
  input  [1:0]  io_in_2_bits_sel_alu3,
  input         io_in_2_bits_mask,
  input  [2:0]  io_in_2_bits_sel_imm,
  input         io_in_2_bits_mem_unsigned,
  input  [5:0]  io_in_2_bits_alu_fn,
  input         io_in_2_bits_mem,
  input  [1:0]  io_in_2_bits_mem_cmd,
  input  [1:0]  io_in_2_bits_mop,
  input  [4:0]  io_in_2_bits_reg_idx1,
  input  [4:0]  io_in_2_bits_reg_idx2,
  input  [4:0]  io_in_2_bits_reg_idx3,
  input  [4:0]  io_in_2_bits_reg_idxw,
  input         io_in_2_bits_wfd,
  input         io_in_2_bits_fence,
  input         io_in_2_bits_sfu,
  input         io_in_2_bits_readmask,
  input         io_in_2_bits_writemask,
  input         io_in_2_bits_wxd,
  input  [31:0] io_in_2_bits_pc,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_inst,
  input  [1:0]  io_in_3_bits_wid,
  input         io_in_3_bits_fp,
  input  [1:0]  io_in_3_bits_branch,
  input         io_in_3_bits_simt_stack,
  input         io_in_3_bits_simt_stack_op,
  input         io_in_3_bits_barrier,
  input  [1:0]  io_in_3_bits_csr,
  input         io_in_3_bits_reverse,
  input  [1:0]  io_in_3_bits_sel_alu2,
  input  [1:0]  io_in_3_bits_sel_alu1,
  input         io_in_3_bits_isvec,
  input  [1:0]  io_in_3_bits_sel_alu3,
  input         io_in_3_bits_mask,
  input  [2:0]  io_in_3_bits_sel_imm,
  input         io_in_3_bits_mem_unsigned,
  input  [5:0]  io_in_3_bits_alu_fn,
  input         io_in_3_bits_mem,
  input  [1:0]  io_in_3_bits_mem_cmd,
  input  [1:0]  io_in_3_bits_mop,
  input  [4:0]  io_in_3_bits_reg_idx1,
  input  [4:0]  io_in_3_bits_reg_idx2,
  input  [4:0]  io_in_3_bits_reg_idx3,
  input  [4:0]  io_in_3_bits_reg_idxw,
  input         io_in_3_bits_wfd,
  input         io_in_3_bits_fence,
  input         io_in_3_bits_sfu,
  input         io_in_3_bits_readmask,
  input         io_in_3_bits_writemask,
  input         io_in_3_bits_wxd,
  input  [31:0] io_in_3_bits_pc,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_inst,
  output [1:0]  io_out_bits_wid,
  output        io_out_bits_fp,
  output [1:0]  io_out_bits_branch,
  output        io_out_bits_simt_stack,
  output        io_out_bits_simt_stack_op,
  output        io_out_bits_barrier,
  output [1:0]  io_out_bits_csr,
  output        io_out_bits_reverse,
  output [1:0]  io_out_bits_sel_alu2,
  output [1:0]  io_out_bits_sel_alu1,
  output        io_out_bits_isvec,
  output [1:0]  io_out_bits_sel_alu3,
  output        io_out_bits_mask,
  output [2:0]  io_out_bits_sel_imm,
  output        io_out_bits_mem_unsigned,
  output [5:0]  io_out_bits_alu_fn,
  output        io_out_bits_mem,
  output [1:0]  io_out_bits_mem_cmd,
  output [1:0]  io_out_bits_mop,
  output [4:0]  io_out_bits_reg_idx1,
  output [4:0]  io_out_bits_reg_idx2,
  output [4:0]  io_out_bits_reg_idx3,
  output [4:0]  io_out_bits_reg_idxw,
  output        io_out_bits_wfd,
  output        io_out_bits_fence,
  output        io_out_bits_sfu,
  output        io_out_bits_readmask,
  output        io_out_bits_writemask,
  output        io_out_bits_wxd,
  output [31:0] io_out_bits_pc
);
  wire  rrarbit_clock; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_ready; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_valid; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_0_bits_inst; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_wid; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_fp; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_branch; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_simt_stack; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_simt_stack_op; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_barrier; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_csr; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_reverse; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_sel_alu2; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_sel_alu1; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_isvec; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_sel_alu3; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_mask; // @[ibuffer.scala 37:21]
  wire [2:0] rrarbit_io_in_0_bits_sel_imm; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_mem_unsigned; // @[ibuffer.scala 37:21]
  wire [5:0] rrarbit_io_in_0_bits_alu_fn; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_mem; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_mem_cmd; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_0_bits_mop; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_0_bits_reg_idx1; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_0_bits_reg_idx2; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_0_bits_reg_idx3; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_0_bits_reg_idxw; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_wfd; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_fence; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_sfu; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_readmask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_writemask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_0_bits_wxd; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_0_bits_pc; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_ready; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_valid; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_1_bits_inst; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_wid; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_fp; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_branch; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_simt_stack; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_simt_stack_op; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_barrier; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_csr; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_reverse; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_sel_alu2; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_sel_alu1; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_isvec; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_sel_alu3; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_mask; // @[ibuffer.scala 37:21]
  wire [2:0] rrarbit_io_in_1_bits_sel_imm; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_mem_unsigned; // @[ibuffer.scala 37:21]
  wire [5:0] rrarbit_io_in_1_bits_alu_fn; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_mem; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_mem_cmd; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_1_bits_mop; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_1_bits_reg_idx1; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_1_bits_reg_idx2; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_1_bits_reg_idx3; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_1_bits_reg_idxw; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_wfd; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_fence; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_sfu; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_readmask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_writemask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_1_bits_wxd; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_1_bits_pc; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_ready; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_valid; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_2_bits_inst; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_wid; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_fp; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_branch; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_simt_stack; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_simt_stack_op; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_barrier; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_csr; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_reverse; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_sel_alu2; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_sel_alu1; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_isvec; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_sel_alu3; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_mask; // @[ibuffer.scala 37:21]
  wire [2:0] rrarbit_io_in_2_bits_sel_imm; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_mem_unsigned; // @[ibuffer.scala 37:21]
  wire [5:0] rrarbit_io_in_2_bits_alu_fn; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_mem; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_mem_cmd; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_2_bits_mop; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_2_bits_reg_idx1; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_2_bits_reg_idx2; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_2_bits_reg_idx3; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_2_bits_reg_idxw; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_wfd; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_fence; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_sfu; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_readmask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_writemask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_2_bits_wxd; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_2_bits_pc; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_ready; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_valid; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_3_bits_inst; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_wid; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_fp; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_branch; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_simt_stack; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_simt_stack_op; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_barrier; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_csr; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_reverse; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_sel_alu2; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_sel_alu1; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_isvec; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_sel_alu3; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_mask; // @[ibuffer.scala 37:21]
  wire [2:0] rrarbit_io_in_3_bits_sel_imm; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_mem_unsigned; // @[ibuffer.scala 37:21]
  wire [5:0] rrarbit_io_in_3_bits_alu_fn; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_mem; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_mem_cmd; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_in_3_bits_mop; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_3_bits_reg_idx1; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_3_bits_reg_idx2; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_3_bits_reg_idx3; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_in_3_bits_reg_idxw; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_wfd; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_fence; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_sfu; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_readmask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_writemask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_in_3_bits_wxd; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_in_3_bits_pc; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_ready; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_valid; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_out_bits_inst; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_wid; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_fp; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_branch; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_simt_stack; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_simt_stack_op; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_barrier; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_csr; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_reverse; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_sel_alu2; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_sel_alu1; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_isvec; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_sel_alu3; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_mask; // @[ibuffer.scala 37:21]
  wire [2:0] rrarbit_io_out_bits_sel_imm; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_mem_unsigned; // @[ibuffer.scala 37:21]
  wire [5:0] rrarbit_io_out_bits_alu_fn; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_mem; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_mem_cmd; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_out_bits_mop; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_out_bits_reg_idx1; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_out_bits_reg_idx2; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_out_bits_reg_idx3; // @[ibuffer.scala 37:21]
  wire [4:0] rrarbit_io_out_bits_reg_idxw; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_wfd; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_fence; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_sfu; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_readmask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_writemask; // @[ibuffer.scala 37:21]
  wire  rrarbit_io_out_bits_wxd; // @[ibuffer.scala 37:21]
  wire [31:0] rrarbit_io_out_bits_pc; // @[ibuffer.scala 37:21]
  wire [1:0] rrarbit_io_chosen; // @[ibuffer.scala 37:21]
  RRArbiter rrarbit ( // @[ibuffer.scala 37:21]
    .clock(rrarbit_clock),
    .io_in_0_ready(rrarbit_io_in_0_ready),
    .io_in_0_valid(rrarbit_io_in_0_valid),
    .io_in_0_bits_inst(rrarbit_io_in_0_bits_inst),
    .io_in_0_bits_wid(rrarbit_io_in_0_bits_wid),
    .io_in_0_bits_fp(rrarbit_io_in_0_bits_fp),
    .io_in_0_bits_branch(rrarbit_io_in_0_bits_branch),
    .io_in_0_bits_simt_stack(rrarbit_io_in_0_bits_simt_stack),
    .io_in_0_bits_simt_stack_op(rrarbit_io_in_0_bits_simt_stack_op),
    .io_in_0_bits_barrier(rrarbit_io_in_0_bits_barrier),
    .io_in_0_bits_csr(rrarbit_io_in_0_bits_csr),
    .io_in_0_bits_reverse(rrarbit_io_in_0_bits_reverse),
    .io_in_0_bits_sel_alu2(rrarbit_io_in_0_bits_sel_alu2),
    .io_in_0_bits_sel_alu1(rrarbit_io_in_0_bits_sel_alu1),
    .io_in_0_bits_isvec(rrarbit_io_in_0_bits_isvec),
    .io_in_0_bits_sel_alu3(rrarbit_io_in_0_bits_sel_alu3),
    .io_in_0_bits_mask(rrarbit_io_in_0_bits_mask),
    .io_in_0_bits_sel_imm(rrarbit_io_in_0_bits_sel_imm),
    .io_in_0_bits_mem_unsigned(rrarbit_io_in_0_bits_mem_unsigned),
    .io_in_0_bits_alu_fn(rrarbit_io_in_0_bits_alu_fn),
    .io_in_0_bits_mem(rrarbit_io_in_0_bits_mem),
    .io_in_0_bits_mem_cmd(rrarbit_io_in_0_bits_mem_cmd),
    .io_in_0_bits_mop(rrarbit_io_in_0_bits_mop),
    .io_in_0_bits_reg_idx1(rrarbit_io_in_0_bits_reg_idx1),
    .io_in_0_bits_reg_idx2(rrarbit_io_in_0_bits_reg_idx2),
    .io_in_0_bits_reg_idx3(rrarbit_io_in_0_bits_reg_idx3),
    .io_in_0_bits_reg_idxw(rrarbit_io_in_0_bits_reg_idxw),
    .io_in_0_bits_wfd(rrarbit_io_in_0_bits_wfd),
    .io_in_0_bits_fence(rrarbit_io_in_0_bits_fence),
    .io_in_0_bits_sfu(rrarbit_io_in_0_bits_sfu),
    .io_in_0_bits_readmask(rrarbit_io_in_0_bits_readmask),
    .io_in_0_bits_writemask(rrarbit_io_in_0_bits_writemask),
    .io_in_0_bits_wxd(rrarbit_io_in_0_bits_wxd),
    .io_in_0_bits_pc(rrarbit_io_in_0_bits_pc),
    .io_in_1_ready(rrarbit_io_in_1_ready),
    .io_in_1_valid(rrarbit_io_in_1_valid),
    .io_in_1_bits_inst(rrarbit_io_in_1_bits_inst),
    .io_in_1_bits_wid(rrarbit_io_in_1_bits_wid),
    .io_in_1_bits_fp(rrarbit_io_in_1_bits_fp),
    .io_in_1_bits_branch(rrarbit_io_in_1_bits_branch),
    .io_in_1_bits_simt_stack(rrarbit_io_in_1_bits_simt_stack),
    .io_in_1_bits_simt_stack_op(rrarbit_io_in_1_bits_simt_stack_op),
    .io_in_1_bits_barrier(rrarbit_io_in_1_bits_barrier),
    .io_in_1_bits_csr(rrarbit_io_in_1_bits_csr),
    .io_in_1_bits_reverse(rrarbit_io_in_1_bits_reverse),
    .io_in_1_bits_sel_alu2(rrarbit_io_in_1_bits_sel_alu2),
    .io_in_1_bits_sel_alu1(rrarbit_io_in_1_bits_sel_alu1),
    .io_in_1_bits_isvec(rrarbit_io_in_1_bits_isvec),
    .io_in_1_bits_sel_alu3(rrarbit_io_in_1_bits_sel_alu3),
    .io_in_1_bits_mask(rrarbit_io_in_1_bits_mask),
    .io_in_1_bits_sel_imm(rrarbit_io_in_1_bits_sel_imm),
    .io_in_1_bits_mem_unsigned(rrarbit_io_in_1_bits_mem_unsigned),
    .io_in_1_bits_alu_fn(rrarbit_io_in_1_bits_alu_fn),
    .io_in_1_bits_mem(rrarbit_io_in_1_bits_mem),
    .io_in_1_bits_mem_cmd(rrarbit_io_in_1_bits_mem_cmd),
    .io_in_1_bits_mop(rrarbit_io_in_1_bits_mop),
    .io_in_1_bits_reg_idx1(rrarbit_io_in_1_bits_reg_idx1),
    .io_in_1_bits_reg_idx2(rrarbit_io_in_1_bits_reg_idx2),
    .io_in_1_bits_reg_idx3(rrarbit_io_in_1_bits_reg_idx3),
    .io_in_1_bits_reg_idxw(rrarbit_io_in_1_bits_reg_idxw),
    .io_in_1_bits_wfd(rrarbit_io_in_1_bits_wfd),
    .io_in_1_bits_fence(rrarbit_io_in_1_bits_fence),
    .io_in_1_bits_sfu(rrarbit_io_in_1_bits_sfu),
    .io_in_1_bits_readmask(rrarbit_io_in_1_bits_readmask),
    .io_in_1_bits_writemask(rrarbit_io_in_1_bits_writemask),
    .io_in_1_bits_wxd(rrarbit_io_in_1_bits_wxd),
    .io_in_1_bits_pc(rrarbit_io_in_1_bits_pc),
    .io_in_2_ready(rrarbit_io_in_2_ready),
    .io_in_2_valid(rrarbit_io_in_2_valid),
    .io_in_2_bits_inst(rrarbit_io_in_2_bits_inst),
    .io_in_2_bits_wid(rrarbit_io_in_2_bits_wid),
    .io_in_2_bits_fp(rrarbit_io_in_2_bits_fp),
    .io_in_2_bits_branch(rrarbit_io_in_2_bits_branch),
    .io_in_2_bits_simt_stack(rrarbit_io_in_2_bits_simt_stack),
    .io_in_2_bits_simt_stack_op(rrarbit_io_in_2_bits_simt_stack_op),
    .io_in_2_bits_barrier(rrarbit_io_in_2_bits_barrier),
    .io_in_2_bits_csr(rrarbit_io_in_2_bits_csr),
    .io_in_2_bits_reverse(rrarbit_io_in_2_bits_reverse),
    .io_in_2_bits_sel_alu2(rrarbit_io_in_2_bits_sel_alu2),
    .io_in_2_bits_sel_alu1(rrarbit_io_in_2_bits_sel_alu1),
    .io_in_2_bits_isvec(rrarbit_io_in_2_bits_isvec),
    .io_in_2_bits_sel_alu3(rrarbit_io_in_2_bits_sel_alu3),
    .io_in_2_bits_mask(rrarbit_io_in_2_bits_mask),
    .io_in_2_bits_sel_imm(rrarbit_io_in_2_bits_sel_imm),
    .io_in_2_bits_mem_unsigned(rrarbit_io_in_2_bits_mem_unsigned),
    .io_in_2_bits_alu_fn(rrarbit_io_in_2_bits_alu_fn),
    .io_in_2_bits_mem(rrarbit_io_in_2_bits_mem),
    .io_in_2_bits_mem_cmd(rrarbit_io_in_2_bits_mem_cmd),
    .io_in_2_bits_mop(rrarbit_io_in_2_bits_mop),
    .io_in_2_bits_reg_idx1(rrarbit_io_in_2_bits_reg_idx1),
    .io_in_2_bits_reg_idx2(rrarbit_io_in_2_bits_reg_idx2),
    .io_in_2_bits_reg_idx3(rrarbit_io_in_2_bits_reg_idx3),
    .io_in_2_bits_reg_idxw(rrarbit_io_in_2_bits_reg_idxw),
    .io_in_2_bits_wfd(rrarbit_io_in_2_bits_wfd),
    .io_in_2_bits_fence(rrarbit_io_in_2_bits_fence),
    .io_in_2_bits_sfu(rrarbit_io_in_2_bits_sfu),
    .io_in_2_bits_readmask(rrarbit_io_in_2_bits_readmask),
    .io_in_2_bits_writemask(rrarbit_io_in_2_bits_writemask),
    .io_in_2_bits_wxd(rrarbit_io_in_2_bits_wxd),
    .io_in_2_bits_pc(rrarbit_io_in_2_bits_pc),
    .io_in_3_ready(rrarbit_io_in_3_ready),
    .io_in_3_valid(rrarbit_io_in_3_valid),
    .io_in_3_bits_inst(rrarbit_io_in_3_bits_inst),
    .io_in_3_bits_wid(rrarbit_io_in_3_bits_wid),
    .io_in_3_bits_fp(rrarbit_io_in_3_bits_fp),
    .io_in_3_bits_branch(rrarbit_io_in_3_bits_branch),
    .io_in_3_bits_simt_stack(rrarbit_io_in_3_bits_simt_stack),
    .io_in_3_bits_simt_stack_op(rrarbit_io_in_3_bits_simt_stack_op),
    .io_in_3_bits_barrier(rrarbit_io_in_3_bits_barrier),
    .io_in_3_bits_csr(rrarbit_io_in_3_bits_csr),
    .io_in_3_bits_reverse(rrarbit_io_in_3_bits_reverse),
    .io_in_3_bits_sel_alu2(rrarbit_io_in_3_bits_sel_alu2),
    .io_in_3_bits_sel_alu1(rrarbit_io_in_3_bits_sel_alu1),
    .io_in_3_bits_isvec(rrarbit_io_in_3_bits_isvec),
    .io_in_3_bits_sel_alu3(rrarbit_io_in_3_bits_sel_alu3),
    .io_in_3_bits_mask(rrarbit_io_in_3_bits_mask),
    .io_in_3_bits_sel_imm(rrarbit_io_in_3_bits_sel_imm),
    .io_in_3_bits_mem_unsigned(rrarbit_io_in_3_bits_mem_unsigned),
    .io_in_3_bits_alu_fn(rrarbit_io_in_3_bits_alu_fn),
    .io_in_3_bits_mem(rrarbit_io_in_3_bits_mem),
    .io_in_3_bits_mem_cmd(rrarbit_io_in_3_bits_mem_cmd),
    .io_in_3_bits_mop(rrarbit_io_in_3_bits_mop),
    .io_in_3_bits_reg_idx1(rrarbit_io_in_3_bits_reg_idx1),
    .io_in_3_bits_reg_idx2(rrarbit_io_in_3_bits_reg_idx2),
    .io_in_3_bits_reg_idx3(rrarbit_io_in_3_bits_reg_idx3),
    .io_in_3_bits_reg_idxw(rrarbit_io_in_3_bits_reg_idxw),
    .io_in_3_bits_wfd(rrarbit_io_in_3_bits_wfd),
    .io_in_3_bits_fence(rrarbit_io_in_3_bits_fence),
    .io_in_3_bits_sfu(rrarbit_io_in_3_bits_sfu),
    .io_in_3_bits_readmask(rrarbit_io_in_3_bits_readmask),
    .io_in_3_bits_writemask(rrarbit_io_in_3_bits_writemask),
    .io_in_3_bits_wxd(rrarbit_io_in_3_bits_wxd),
    .io_in_3_bits_pc(rrarbit_io_in_3_bits_pc),
    .io_out_ready(rrarbit_io_out_ready),
    .io_out_valid(rrarbit_io_out_valid),
    .io_out_bits_inst(rrarbit_io_out_bits_inst),
    .io_out_bits_wid(rrarbit_io_out_bits_wid),
    .io_out_bits_fp(rrarbit_io_out_bits_fp),
    .io_out_bits_branch(rrarbit_io_out_bits_branch),
    .io_out_bits_simt_stack(rrarbit_io_out_bits_simt_stack),
    .io_out_bits_simt_stack_op(rrarbit_io_out_bits_simt_stack_op),
    .io_out_bits_barrier(rrarbit_io_out_bits_barrier),
    .io_out_bits_csr(rrarbit_io_out_bits_csr),
    .io_out_bits_reverse(rrarbit_io_out_bits_reverse),
    .io_out_bits_sel_alu2(rrarbit_io_out_bits_sel_alu2),
    .io_out_bits_sel_alu1(rrarbit_io_out_bits_sel_alu1),
    .io_out_bits_isvec(rrarbit_io_out_bits_isvec),
    .io_out_bits_sel_alu3(rrarbit_io_out_bits_sel_alu3),
    .io_out_bits_mask(rrarbit_io_out_bits_mask),
    .io_out_bits_sel_imm(rrarbit_io_out_bits_sel_imm),
    .io_out_bits_mem_unsigned(rrarbit_io_out_bits_mem_unsigned),
    .io_out_bits_alu_fn(rrarbit_io_out_bits_alu_fn),
    .io_out_bits_mem(rrarbit_io_out_bits_mem),
    .io_out_bits_mem_cmd(rrarbit_io_out_bits_mem_cmd),
    .io_out_bits_mop(rrarbit_io_out_bits_mop),
    .io_out_bits_reg_idx1(rrarbit_io_out_bits_reg_idx1),
    .io_out_bits_reg_idx2(rrarbit_io_out_bits_reg_idx2),
    .io_out_bits_reg_idx3(rrarbit_io_out_bits_reg_idx3),
    .io_out_bits_reg_idxw(rrarbit_io_out_bits_reg_idxw),
    .io_out_bits_wfd(rrarbit_io_out_bits_wfd),
    .io_out_bits_fence(rrarbit_io_out_bits_fence),
    .io_out_bits_sfu(rrarbit_io_out_bits_sfu),
    .io_out_bits_readmask(rrarbit_io_out_bits_readmask),
    .io_out_bits_writemask(rrarbit_io_out_bits_writemask),
    .io_out_bits_wxd(rrarbit_io_out_bits_wxd),
    .io_out_bits_pc(rrarbit_io_out_bits_pc),
    .io_chosen(rrarbit_io_chosen)
  );
  assign io_in_0_ready = rrarbit_io_in_0_ready; // @[ibuffer.scala 38:16]
  assign io_in_1_ready = rrarbit_io_in_1_ready; // @[ibuffer.scala 38:16]
  assign io_in_2_ready = rrarbit_io_in_2_ready; // @[ibuffer.scala 38:16]
  assign io_in_3_ready = rrarbit_io_in_3_ready; // @[ibuffer.scala 38:16]
  assign io_out_valid = rrarbit_io_out_valid; // @[ibuffer.scala 39:9]
  assign io_out_bits_inst = rrarbit_io_out_bits_inst; // @[ibuffer.scala 39:9]
  assign io_out_bits_wid = rrarbit_io_out_bits_wid; // @[ibuffer.scala 39:9]
  assign io_out_bits_fp = rrarbit_io_out_bits_fp; // @[ibuffer.scala 39:9]
  assign io_out_bits_branch = rrarbit_io_out_bits_branch; // @[ibuffer.scala 39:9]
  assign io_out_bits_simt_stack = rrarbit_io_out_bits_simt_stack; // @[ibuffer.scala 39:9]
  assign io_out_bits_simt_stack_op = rrarbit_io_out_bits_simt_stack_op; // @[ibuffer.scala 39:9]
  assign io_out_bits_barrier = rrarbit_io_out_bits_barrier; // @[ibuffer.scala 39:9]
  assign io_out_bits_csr = rrarbit_io_out_bits_csr; // @[ibuffer.scala 39:9]
  assign io_out_bits_reverse = rrarbit_io_out_bits_reverse; // @[ibuffer.scala 39:9]
  assign io_out_bits_sel_alu2 = rrarbit_io_out_bits_sel_alu2; // @[ibuffer.scala 39:9]
  assign io_out_bits_sel_alu1 = rrarbit_io_out_bits_sel_alu1; // @[ibuffer.scala 39:9]
  assign io_out_bits_isvec = rrarbit_io_out_bits_isvec; // @[ibuffer.scala 39:9]
  assign io_out_bits_sel_alu3 = rrarbit_io_out_bits_sel_alu3; // @[ibuffer.scala 39:9]
  assign io_out_bits_mask = rrarbit_io_out_bits_mask; // @[ibuffer.scala 39:9]
  assign io_out_bits_sel_imm = rrarbit_io_out_bits_sel_imm; // @[ibuffer.scala 39:9]
  assign io_out_bits_mem_unsigned = rrarbit_io_out_bits_mem_unsigned; // @[ibuffer.scala 39:9]
  assign io_out_bits_alu_fn = rrarbit_io_out_bits_alu_fn; // @[ibuffer.scala 39:9]
  assign io_out_bits_mem = rrarbit_io_out_bits_mem; // @[ibuffer.scala 39:9]
  assign io_out_bits_mem_cmd = rrarbit_io_out_bits_mem_cmd; // @[ibuffer.scala 39:9]
  assign io_out_bits_mop = rrarbit_io_out_bits_mop; // @[ibuffer.scala 39:9]
  assign io_out_bits_reg_idx1 = rrarbit_io_out_bits_reg_idx1; // @[ibuffer.scala 39:9]
  assign io_out_bits_reg_idx2 = rrarbit_io_out_bits_reg_idx2; // @[ibuffer.scala 39:9]
  assign io_out_bits_reg_idx3 = rrarbit_io_out_bits_reg_idx3; // @[ibuffer.scala 39:9]
  assign io_out_bits_reg_idxw = rrarbit_io_out_bits_reg_idxw; // @[ibuffer.scala 39:9]
  assign io_out_bits_wfd = rrarbit_io_out_bits_wfd; // @[ibuffer.scala 39:9]
  assign io_out_bits_fence = rrarbit_io_out_bits_fence; // @[ibuffer.scala 39:9]
  assign io_out_bits_sfu = rrarbit_io_out_bits_sfu; // @[ibuffer.scala 39:9]
  assign io_out_bits_readmask = rrarbit_io_out_bits_readmask; // @[ibuffer.scala 39:9]
  assign io_out_bits_writemask = rrarbit_io_out_bits_writemask; // @[ibuffer.scala 39:9]
  assign io_out_bits_wxd = rrarbit_io_out_bits_wxd; // @[ibuffer.scala 39:9]
  assign io_out_bits_pc = rrarbit_io_out_bits_pc; // @[ibuffer.scala 39:9]
  assign rrarbit_clock = clock;
  assign rrarbit_io_in_0_valid = io_in_0_valid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_inst = io_in_0_bits_inst; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_wid = io_in_0_bits_wid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_fp = io_in_0_bits_fp; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_branch = io_in_0_bits_branch; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_simt_stack = io_in_0_bits_simt_stack; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_simt_stack_op = io_in_0_bits_simt_stack_op; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_barrier = io_in_0_bits_barrier; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_csr = io_in_0_bits_csr; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_reverse = io_in_0_bits_reverse; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_sel_alu2 = io_in_0_bits_sel_alu2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_sel_alu1 = io_in_0_bits_sel_alu1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_isvec = io_in_0_bits_isvec; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_sel_alu3 = io_in_0_bits_sel_alu3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_mask = io_in_0_bits_mask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_sel_imm = io_in_0_bits_sel_imm; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_mem_unsigned = io_in_0_bits_mem_unsigned; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_alu_fn = io_in_0_bits_alu_fn; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_mem = io_in_0_bits_mem; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_mem_cmd = io_in_0_bits_mem_cmd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_mop = io_in_0_bits_mop; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_reg_idx1 = io_in_0_bits_reg_idx1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_reg_idx2 = io_in_0_bits_reg_idx2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_reg_idx3 = io_in_0_bits_reg_idx3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_reg_idxw = io_in_0_bits_reg_idxw; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_wfd = io_in_0_bits_wfd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_fence = io_in_0_bits_fence; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_sfu = io_in_0_bits_sfu; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_readmask = io_in_0_bits_readmask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_writemask = io_in_0_bits_writemask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_wxd = io_in_0_bits_wxd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_0_bits_pc = io_in_0_bits_pc; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_valid = io_in_1_valid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_inst = io_in_1_bits_inst; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_wid = io_in_1_bits_wid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_fp = io_in_1_bits_fp; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_branch = io_in_1_bits_branch; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_simt_stack = io_in_1_bits_simt_stack; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_simt_stack_op = io_in_1_bits_simt_stack_op; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_barrier = io_in_1_bits_barrier; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_csr = io_in_1_bits_csr; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_reverse = io_in_1_bits_reverse; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_sel_alu2 = io_in_1_bits_sel_alu2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_sel_alu1 = io_in_1_bits_sel_alu1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_isvec = io_in_1_bits_isvec; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_sel_alu3 = io_in_1_bits_sel_alu3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_mask = io_in_1_bits_mask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_sel_imm = io_in_1_bits_sel_imm; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_mem_unsigned = io_in_1_bits_mem_unsigned; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_alu_fn = io_in_1_bits_alu_fn; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_mem = io_in_1_bits_mem; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_mem_cmd = io_in_1_bits_mem_cmd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_mop = io_in_1_bits_mop; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_reg_idx1 = io_in_1_bits_reg_idx1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_reg_idx2 = io_in_1_bits_reg_idx2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_reg_idx3 = io_in_1_bits_reg_idx3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_reg_idxw = io_in_1_bits_reg_idxw; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_wfd = io_in_1_bits_wfd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_fence = io_in_1_bits_fence; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_sfu = io_in_1_bits_sfu; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_readmask = io_in_1_bits_readmask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_writemask = io_in_1_bits_writemask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_wxd = io_in_1_bits_wxd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_1_bits_pc = io_in_1_bits_pc; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_valid = io_in_2_valid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_inst = io_in_2_bits_inst; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_wid = io_in_2_bits_wid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_fp = io_in_2_bits_fp; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_branch = io_in_2_bits_branch; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_simt_stack = io_in_2_bits_simt_stack; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_simt_stack_op = io_in_2_bits_simt_stack_op; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_barrier = io_in_2_bits_barrier; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_csr = io_in_2_bits_csr; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_reverse = io_in_2_bits_reverse; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_sel_alu2 = io_in_2_bits_sel_alu2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_sel_alu1 = io_in_2_bits_sel_alu1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_isvec = io_in_2_bits_isvec; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_sel_alu3 = io_in_2_bits_sel_alu3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_mask = io_in_2_bits_mask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_sel_imm = io_in_2_bits_sel_imm; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_mem_unsigned = io_in_2_bits_mem_unsigned; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_alu_fn = io_in_2_bits_alu_fn; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_mem = io_in_2_bits_mem; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_mem_cmd = io_in_2_bits_mem_cmd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_mop = io_in_2_bits_mop; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_reg_idx1 = io_in_2_bits_reg_idx1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_reg_idx2 = io_in_2_bits_reg_idx2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_reg_idx3 = io_in_2_bits_reg_idx3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_reg_idxw = io_in_2_bits_reg_idxw; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_wfd = io_in_2_bits_wfd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_fence = io_in_2_bits_fence; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_sfu = io_in_2_bits_sfu; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_readmask = io_in_2_bits_readmask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_writemask = io_in_2_bits_writemask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_wxd = io_in_2_bits_wxd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_2_bits_pc = io_in_2_bits_pc; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_valid = io_in_3_valid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_inst = io_in_3_bits_inst; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_wid = io_in_3_bits_wid; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_fp = io_in_3_bits_fp; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_branch = io_in_3_bits_branch; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_simt_stack = io_in_3_bits_simt_stack; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_simt_stack_op = io_in_3_bits_simt_stack_op; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_barrier = io_in_3_bits_barrier; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_csr = io_in_3_bits_csr; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_reverse = io_in_3_bits_reverse; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_sel_alu2 = io_in_3_bits_sel_alu2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_sel_alu1 = io_in_3_bits_sel_alu1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_isvec = io_in_3_bits_isvec; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_sel_alu3 = io_in_3_bits_sel_alu3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_mask = io_in_3_bits_mask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_sel_imm = io_in_3_bits_sel_imm; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_mem_unsigned = io_in_3_bits_mem_unsigned; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_alu_fn = io_in_3_bits_alu_fn; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_mem = io_in_3_bits_mem; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_mem_cmd = io_in_3_bits_mem_cmd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_mop = io_in_3_bits_mop; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_reg_idx1 = io_in_3_bits_reg_idx1; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_reg_idx2 = io_in_3_bits_reg_idx2; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_reg_idx3 = io_in_3_bits_reg_idx3; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_reg_idxw = io_in_3_bits_reg_idxw; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_wfd = io_in_3_bits_wfd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_fence = io_in_3_bits_fence; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_sfu = io_in_3_bits_sfu; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_readmask = io_in_3_bits_readmask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_writemask = io_in_3_bits_writemask; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_wxd = io_in_3_bits_wxd; // @[ibuffer.scala 38:16]
  assign rrarbit_io_in_3_bits_pc = io_in_3_bits_pc; // @[ibuffer.scala 38:16]
  assign rrarbit_io_out_ready = io_out_ready; // @[ibuffer.scala 39:9]
endmodule
module Queue_46(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_wid,
  input  [31:0] io_enq_bits_PC_branch,
  input  [7:0]  io_enq_bits_mask_init,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_opcode,
  output [1:0]  io_deq_bits_wid,
  output [31:0] io_deq_bits_PC_branch,
  output [7:0]  io_deq_bits_mask_init
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_opcode [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_PC_branch [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_PC_branch_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_PC_branch_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_PC_branch_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_PC_branch_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_PC_branch_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_PC_branch_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_PC_branch_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask_init [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_init_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_init_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_init_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_init_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_init_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_init_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_init_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wid_io_deq_bits_MPORT_data = ram_wid[ram_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wid_MPORT_data = io_enq_bits_wid;
  assign ram_wid_MPORT_addr = 1'h0;
  assign ram_wid_MPORT_mask = 1'h1;
  assign ram_wid_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_PC_branch_io_deq_bits_MPORT_en = 1'h1;
  assign ram_PC_branch_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_PC_branch_io_deq_bits_MPORT_data = ram_PC_branch[ram_PC_branch_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_PC_branch_MPORT_data = io_enq_bits_PC_branch;
  assign ram_PC_branch_MPORT_addr = 1'h0;
  assign ram_PC_branch_MPORT_mask = 1'h1;
  assign ram_PC_branch_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_mask_init_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_init_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_init_io_deq_bits_MPORT_data = ram_mask_init[ram_mask_init_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_init_MPORT_data = io_enq_bits_mask_init;
  assign ram_mask_init_MPORT_addr = 1'h0;
  assign ram_mask_init_MPORT_mask = 1'h1;
  assign ram_mask_init_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_opcode = empty ? io_enq_bits_opcode : ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_wid = empty ? io_enq_bits_wid : ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_PC_branch = empty ? io_enq_bits_PC_branch : ram_PC_branch_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_mask_init = empty ? io_enq_bits_mask_init : ram_mask_init_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wid_MPORT_en & ram_wid_MPORT_mask) begin
      ram_wid[ram_wid_MPORT_addr] <= ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_PC_branch_MPORT_en & ram_PC_branch_MPORT_mask) begin
      ram_PC_branch[ram_PC_branch_MPORT_addr] <= ram_PC_branch_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_init_MPORT_en & ram_mask_init_MPORT_mask) begin
      ram_mask_init[ram_mask_init_MPORT_addr] <= ram_mask_init_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wid[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_PC_branch[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask_init[initvar] = _RAND_3[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_47(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_wid,
  input         io_enq_bits_jump,
  input  [31:0] io_enq_bits_new_pc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_wid,
  output        io_deq_bits_jump,
  output [31:0] io_deq_bits_new_pc
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_wid [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wid_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_jump [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_jump_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_jump_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_jump_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_jump_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_new_pc [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_new_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_new_pc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_new_pc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_11 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_11 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  assign ram_wid_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wid_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wid_io_deq_bits_MPORT_data = ram_wid[ram_wid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wid_MPORT_data = io_enq_bits_wid;
  assign ram_wid_MPORT_addr = 1'h0;
  assign ram_wid_MPORT_mask = 1'h1;
  assign ram_wid_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_jump_io_deq_bits_MPORT_en = 1'h1;
  assign ram_jump_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_jump_io_deq_bits_MPORT_data = ram_jump[ram_jump_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_jump_MPORT_data = io_enq_bits_jump;
  assign ram_jump_MPORT_addr = 1'h0;
  assign ram_jump_MPORT_mask = 1'h1;
  assign ram_jump_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_new_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_new_pc_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_new_pc_io_deq_bits_MPORT_data = ram_new_pc[ram_new_pc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_new_pc_MPORT_data = io_enq_bits_new_pc;
  assign ram_new_pc_MPORT_addr = 1'h0;
  assign ram_new_pc_MPORT_mask = 1'h1;
  assign ram_new_pc_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_wid = empty ? io_enq_bits_wid : ram_wid_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_jump = empty ? io_enq_bits_jump : ram_jump_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_new_pc = empty ? io_enq_bits_new_pc : ram_new_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  always @(posedge clock) begin
    if (ram_wid_MPORT_en & ram_wid_MPORT_mask) begin
      ram_wid[ram_wid_MPORT_addr] <= ram_wid_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_jump_MPORT_en & ram_jump_MPORT_mask) begin
      ram_jump[ram_jump_MPORT_addr] <= ram_jump_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_new_pc_MPORT_en & ram_new_pc_MPORT_mask) begin
      ram_new_pc[ram_new_pc_MPORT_addr] <= ram_new_pc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      if (empty) begin // @[Decoupled.scala 301:17]
        if (io_deq_ready) begin // @[Decoupled.scala 304:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 304:35]
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wid[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_jump[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_new_pc[initvar] = _RAND_2[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ipdom_stack(
  input         clock,
  input         reset,
  input         io_push,
  input         io_pop,
  input         io_pair,
  input         io_branchImm,
  input  [39:0] io_q1,
  input  [39:0] io_q2,
  output [39:0] io_d,
  output        io_index,
  output        io_pairo
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [79:0] stack_mem [0:7]; // @[SIMT_STACK.scala 40:22]
  wire  stack_mem_dout_MPORT_en; // @[SIMT_STACK.scala 40:22]
  wire [2:0] stack_mem_dout_MPORT_addr; // @[SIMT_STACK.scala 40:22]
  wire [79:0] stack_mem_dout_MPORT_data; // @[SIMT_STACK.scala 40:22]
  wire [79:0] stack_mem_MPORT_data; // @[SIMT_STACK.scala 40:22]
  wire [2:0] stack_mem_MPORT_addr; // @[SIMT_STACK.scala 40:22]
  wire  stack_mem_MPORT_mask; // @[SIMT_STACK.scala 40:22]
  wire  stack_mem_MPORT_en; // @[SIMT_STACK.scala 40:22]
  reg  is_part_0; // @[SIMT_STACK.scala 36:24]
  reg  is_part_1; // @[SIMT_STACK.scala 36:24]
  reg  is_part_2; // @[SIMT_STACK.scala 36:24]
  reg  is_part_3; // @[SIMT_STACK.scala 36:24]
  reg  is_part_4; // @[SIMT_STACK.scala 36:24]
  reg  is_part_5; // @[SIMT_STACK.scala 36:24]
  reg  is_part_6; // @[SIMT_STACK.scala 36:24]
  reg  is_part_7; // @[SIMT_STACK.scala 36:24]
  reg [3:0] rd_ptr; // @[SIMT_STACK.scala 37:24]
  reg [3:0] wr_ptr; // @[SIMT_STACK.scala 38:24]
  reg  pair_mem_0; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_1; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_2; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_3; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_4; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_5; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_6; // @[SIMT_STACK.scala 42:25]
  reg  pair_mem_7; // @[SIMT_STACK.scala 42:25]
  wire  diverge = ~io_pair | io_branchImm; // @[SIMT_STACK.scala 50:23]
  wire [3:0] _wr_ptr_T_1 = wr_ptr + 4'h1; // @[SIMT_STACK.scala 54:23]
  wire  _GEN_8 = 3'h0 == wr_ptr[2:0] ? io_pair : pair_mem_0; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_9 = 3'h1 == wr_ptr[2:0] ? io_pair : pair_mem_1; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_10 = 3'h2 == wr_ptr[2:0] ? io_pair : pair_mem_2; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_11 = 3'h3 == wr_ptr[2:0] ? io_pair : pair_mem_3; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_12 = 3'h4 == wr_ptr[2:0] ? io_pair : pair_mem_4; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_13 = 3'h5 == wr_ptr[2:0] ? io_pair : pair_mem_5; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_14 = 3'h6 == wr_ptr[2:0] ? io_pair : pair_mem_6; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_15 = 3'h7 == wr_ptr[2:0] ? io_pair : pair_mem_7; // @[SIMT_STACK.scala 56:{22,22} 42:25]
  wire  _GEN_17 = 3'h1 == rd_ptr[2:0] ? is_part_1 : is_part_0; // @[SIMT_STACK.scala 61:{23,23}]
  wire  _GEN_18 = 3'h2 == rd_ptr[2:0] ? is_part_2 : _GEN_17; // @[SIMT_STACK.scala 61:{23,23}]
  wire  _GEN_19 = 3'h3 == rd_ptr[2:0] ? is_part_3 : _GEN_18; // @[SIMT_STACK.scala 61:{23,23}]
  wire  _GEN_20 = 3'h4 == rd_ptr[2:0] ? is_part_4 : _GEN_19; // @[SIMT_STACK.scala 61:{23,23}]
  wire  _GEN_21 = 3'h5 == rd_ptr[2:0] ? is_part_5 : _GEN_20; // @[SIMT_STACK.scala 61:{23,23}]
  wire  _GEN_22 = 3'h6 == rd_ptr[2:0] ? is_part_6 : _GEN_21; // @[SIMT_STACK.scala 61:{23,23}]
  wire  _GEN_23 = 3'h7 == rd_ptr[2:0] ? is_part_7 : _GEN_22; // @[SIMT_STACK.scala 61:{23,23}]
  wire [3:0] _GEN_91 = {{3'd0}, _GEN_23}; // @[SIMT_STACK.scala 61:23]
  wire [3:0] _wr_ptr_T_4 = wr_ptr - _GEN_91; // @[SIMT_STACK.scala 61:23]
  wire [3:0] _rd_ptr_T_2 = rd_ptr - _GEN_91; // @[SIMT_STACK.scala 62:23]
  wire  _GEN_32 = 3'h0 == rd_ptr[2:0] | is_part_0; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_33 = 3'h1 == rd_ptr[2:0] | is_part_1; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_34 = 3'h2 == rd_ptr[2:0] | is_part_2; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_35 = 3'h3 == rd_ptr[2:0] | is_part_3; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_36 = 3'h4 == rd_ptr[2:0] | is_part_4; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_37 = 3'h5 == rd_ptr[2:0] | is_part_5; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_38 = 3'h6 == rd_ptr[2:0] | is_part_6; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_39 = 3'h7 == rd_ptr[2:0] | is_part_7; // @[SIMT_STACK.scala 63:{21,21} 36:24]
  wire  _GEN_60 = io_push ? _GEN_8 : pair_mem_0; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_61 = io_push ? _GEN_9 : pair_mem_1; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_62 = io_push ? _GEN_10 : pair_mem_2; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_63 = io_push ? _GEN_11 : pair_mem_3; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_64 = io_push ? _GEN_12 : pair_mem_4; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_65 = io_push ? _GEN_13 : pair_mem_5; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_66 = io_push ? _GEN_14 : pair_mem_6; // @[SIMT_STACK.scala 52:17 42:25]
  wire  _GEN_67 = io_push ? _GEN_15 : pair_mem_7; // @[SIMT_STACK.scala 52:17 42:25]
  wire [79:0] dout = stack_mem_dout_MPORT_data;
  wire [40:0] _io_d_T_2 = io_index ? {{1'd0}, dout[79:40]} : dout[40:0]; // @[SIMT_STACK.scala 69:18]
  wire  _GEN_82 = 3'h1 == rd_ptr[2:0] ? pair_mem_1 : pair_mem_0; // @[SIMT_STACK.scala 71:{12,12}]
  wire  _GEN_83 = 3'h2 == rd_ptr[2:0] ? pair_mem_2 : _GEN_82; // @[SIMT_STACK.scala 71:{12,12}]
  wire  _GEN_84 = 3'h3 == rd_ptr[2:0] ? pair_mem_3 : _GEN_83; // @[SIMT_STACK.scala 71:{12,12}]
  wire  _GEN_85 = 3'h4 == rd_ptr[2:0] ? pair_mem_4 : _GEN_84; // @[SIMT_STACK.scala 71:{12,12}]
  wire  _GEN_86 = 3'h5 == rd_ptr[2:0] ? pair_mem_5 : _GEN_85; // @[SIMT_STACK.scala 71:{12,12}]
  wire  _GEN_87 = 3'h6 == rd_ptr[2:0] ? pair_mem_6 : _GEN_86; // @[SIMT_STACK.scala 71:{12,12}]
  assign stack_mem_dout_MPORT_en = 1'h1;
  assign stack_mem_dout_MPORT_addr = rd_ptr[2:0];
  assign stack_mem_dout_MPORT_data = stack_mem[stack_mem_dout_MPORT_addr]; // @[SIMT_STACK.scala 40:22]
  assign stack_mem_MPORT_data = {io_q1,io_q2};
  assign stack_mem_MPORT_addr = wr_ptr[2:0];
  assign stack_mem_MPORT_mask = 1'h1;
  assign stack_mem_MPORT_en = io_push;
  assign io_d = _io_d_T_2[39:0]; // @[SIMT_STACK.scala 69:12]
  assign io_index = 3'h7 == rd_ptr[2:0] ? is_part_7 : _GEN_22; // @[SIMT_STACK.scala 68:{37,37}]
  assign io_pairo = 3'h7 == rd_ptr[2:0] ? pair_mem_7 : _GEN_87; // @[SIMT_STACK.scala 71:{12,12}]
  always @(posedge clock) begin
    if (stack_mem_MPORT_en & stack_mem_MPORT_mask) begin
      stack_mem[stack_mem_MPORT_addr] <= stack_mem_MPORT_data; // @[SIMT_STACK.scala 40:22]
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_0 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h0 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_0 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_0 <= _GEN_32;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_1 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h1 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_1 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_1 <= _GEN_33;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_2 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h2 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_2 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_2 <= _GEN_34;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_3 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h3 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_3 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_3 <= _GEN_35;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_4 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h4 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_4 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_4 <= _GEN_36;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_5 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h5 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_5 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_5 <= _GEN_37;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_6 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h6 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_6 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_6 <= _GEN_38;
    end
    if (reset) begin // @[SIMT_STACK.scala 36:24]
      is_part_7 <= 1'h0; // @[SIMT_STACK.scala 36:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      if (3'h7 == wr_ptr[2:0]) begin // @[SIMT_STACK.scala 55:21]
        is_part_7 <= diverge; // @[SIMT_STACK.scala 55:21]
      end
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      is_part_7 <= _GEN_39;
    end
    if (reset) begin // @[SIMT_STACK.scala 37:24]
      rd_ptr <= 4'h0; // @[SIMT_STACK.scala 37:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      rd_ptr <= wr_ptr; // @[SIMT_STACK.scala 53:13]
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      rd_ptr <= _rd_ptr_T_2; // @[SIMT_STACK.scala 62:13]
    end
    if (reset) begin // @[SIMT_STACK.scala 38:24]
      wr_ptr <= 4'h0; // @[SIMT_STACK.scala 38:24]
    end else if (io_push) begin // @[SIMT_STACK.scala 52:17]
      wr_ptr <= _wr_ptr_T_1; // @[SIMT_STACK.scala 54:13]
    end else if (io_pop) begin // @[SIMT_STACK.scala 60:23]
      wr_ptr <= _wr_ptr_T_4; // @[SIMT_STACK.scala 61:13]
    end
    pair_mem_0 <= reset | _GEN_60; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_1 <= reset | _GEN_61; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_2 <= reset | _GEN_62; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_3 <= reset | _GEN_63; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_4 <= reset | _GEN_64; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_5 <= reset | _GEN_65; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_6 <= reset | _GEN_66; // @[SIMT_STACK.scala 42:{25,25}]
    pair_mem_7 <= reset | _GEN_67; // @[SIMT_STACK.scala 42:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    stack_mem[initvar] = _RAND_0[79:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  is_part_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  is_part_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  is_part_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  is_part_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  is_part_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  is_part_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  is_part_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  is_part_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rd_ptr = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  wr_ptr = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  pair_mem_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pair_mem_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  pair_mem_2 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pair_mem_3 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  pair_mem_4 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pair_mem_5 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  pair_mem_6 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pair_mem_7 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SIMT_STACK(
  input         clock,
  input         reset,
  output        io_branch_ctl_ready,
  input         io_branch_ctl_valid,
  input         io_branch_ctl_bits_opcode,
  input  [1:0]  io_branch_ctl_bits_wid,
  input  [31:0] io_branch_ctl_bits_PC_branch,
  input  [7:0]  io_branch_ctl_bits_mask_init,
  output        io_if_mask_ready,
  input         io_if_mask_valid,
  input  [7:0]  io_if_mask_bits_if_mask,
  input  [1:0]  io_if_mask_bits_wid,
  input  [1:0]  io_input_wid,
  output [7:0]  io_out_mask,
  output        io_complete_valid,
  output [1:0]  io_complete_bits,
  input         io_fetch_ctl_ready,
  output        io_fetch_ctl_valid,
  output [1:0]  io_fetch_ctl_bits_wid,
  output        io_fetch_ctl_bits_jump,
  output [31:0] io_fetch_ctl_bits_new_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  branch_ctl_buf_clock; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_reset; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [1:0] branch_ctl_buf_io_enq_bits_wid; // @[Decoupled.scala 361:21]
  wire [31:0] branch_ctl_buf_io_enq_bits_PC_branch; // @[Decoupled.scala 361:21]
  wire [7:0] branch_ctl_buf_io_enq_bits_mask_init; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  branch_ctl_buf_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [1:0] branch_ctl_buf_io_deq_bits_wid; // @[Decoupled.scala 361:21]
  wire [31:0] branch_ctl_buf_io_deq_bits_PC_branch; // @[Decoupled.scala 361:21]
  wire [7:0] branch_ctl_buf_io_deq_bits_mask_init; // @[Decoupled.scala 361:21]
  wire  fetch_ctl_buf_clock; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_reset; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_io_enq_ready; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_io_enq_valid; // @[SIMT_STACK.scala 133:29]
  wire [1:0] fetch_ctl_buf_io_enq_bits_wid; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_io_enq_bits_jump; // @[SIMT_STACK.scala 133:29]
  wire [31:0] fetch_ctl_buf_io_enq_bits_new_pc; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_io_deq_ready; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_io_deq_valid; // @[SIMT_STACK.scala 133:29]
  wire [1:0] fetch_ctl_buf_io_deq_bits_wid; // @[SIMT_STACK.scala 133:29]
  wire  fetch_ctl_buf_io_deq_bits_jump; // @[SIMT_STACK.scala 133:29]
  wire [31:0] fetch_ctl_buf_io_deq_bits_new_pc; // @[SIMT_STACK.scala 133:29]
  wire  ipdom_stack_clock; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_reset; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_io_push; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_io_pop; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_io_pair; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_io_branchImm; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_io_q1; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_io_q2; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_io_d; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_io_index; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_io_pairo; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_clock; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_reset; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_io_push; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_io_pop; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_io_pair; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_io_branchImm; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_1_io_q1; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_1_io_q2; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_1_io_d; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_io_index; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_1_io_pairo; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_clock; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_reset; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_io_push; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_io_pop; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_io_pair; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_io_branchImm; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_2_io_q1; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_2_io_q2; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_2_io_d; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_io_index; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_2_io_pairo; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_clock; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_reset; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_io_push; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_io_pop; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_io_pair; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_io_branchImm; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_3_io_q1; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_3_io_q2; // @[SIMT_STACK.scala 160:55]
  wire [39:0] ipdom_stack_3_io_d; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_io_index; // @[SIMT_STACK.scala 160:55]
  wire  ipdom_stack_3_io_pairo; // @[SIMT_STACK.scala 160:55]
  reg [7:0] thread_masks_0; // @[SIMT_STACK.scala 137:29]
  reg [7:0] thread_masks_1; // @[SIMT_STACK.scala 137:29]
  reg [7:0] thread_masks_2; // @[SIMT_STACK.scala 137:29]
  reg [7:0] thread_masks_3; // @[SIMT_STACK.scala 137:29]
  wire  opcode = branch_ctl_buf_io_deq_bits_opcode; // @[SIMT_STACK.scala 123:26 162:10]
  wire  _T = ~opcode; // @[SIMT_STACK.scala 166:39]
  wire  if_mask_buf_ready = fetch_ctl_buf_io_enq_ready; // @[Decoupled.scala 355:21 SIMT_STACK.scala 195:21]
  wire  _branch_ctl_buf_io_deq_ready_T = if_mask_buf_ready & io_if_mask_valid; // @[Decoupled.scala 50:35]
  wire  _T_5 = branch_ctl_buf_io_deq_valid & opcode; // @[SIMT_STACK.scala 179:35]
  wire  _GEN_1 = branch_ctl_buf_io_deq_valid & ~opcode & branch_ctl_buf_io_deq_bits_wid == io_if_mask_bits_wid ?
    _branch_ctl_buf_io_deq_ready_T : _T_5; // @[SIMT_STACK.scala 166:102 167:26]
  wire [7:0] if_mask = io_if_mask_bits_if_mask & branch_ctl_buf_io_deq_bits_mask_init; // @[SIMT_STACK.scala 186:40]
  wire [7:0] _else_mask_T = ~io_if_mask_bits_if_mask; // @[SIMT_STACK.scala 187:16]
  wire [7:0] else_mask = _else_mask_T & branch_ctl_buf_io_deq_bits_mask_init; // @[SIMT_STACK.scala 187:51]
  wire [1:0] warp_id = branch_ctl_buf_io_deq_bits_wid; // @[SIMT_STACK.scala 124:26 164:12]
  wire [7:0] _GEN_4 = 2'h1 == warp_id ? thread_masks_1 : thread_masks_0; // @[SIMT_STACK.scala 191:{26,26}]
  wire [7:0] _GEN_5 = 2'h2 == warp_id ? thread_masks_2 : _GEN_4; // @[SIMT_STACK.scala 191:{26,26}]
  wire [7:0] _GEN_6 = 2'h3 == warp_id ? thread_masks_3 : _GEN_5; // @[SIMT_STACK.scala 191:{26,26}]
  wire [7:0] _diverge_T = else_mask & _GEN_6; // @[SIMT_STACK.scala 192:27]
  wire  elseOnly = _branch_ctl_buf_io_deq_ready_T & else_mask == _GEN_6; // @[SIMT_STACK.scala 189:12 190:28 191:13]
  wire  _io_complete_valid_T_4 = ~elseOnly; // @[SIMT_STACK.scala 196:77]
  wire  _push_0_T_1 = branch_ctl_buf_io_deq_ready & branch_ctl_buf_io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _push_0_T_3 = 2'h0 == warp_id; // @[SIMT_STACK.scala 200:75]
  wire [31:0] PC_branch = branch_ctl_buf_io_deq_bits_PC_branch; // @[SIMT_STACK.scala 125:26 163:13]
  wire  ipdom_stack_4_0_index = ipdom_stack_io_index; // @[SIMT_STACK.scala 160:{29,29}]
  wire  ipdom_index_0 = ~ipdom_stack_4_0_index; // @[SIMT_STACK.scala 229:28]
  wire  _push_1_T_3 = 2'h1 == warp_id; // @[SIMT_STACK.scala 200:75]
  wire  ipdom_stack_4_1_index = ipdom_stack_1_io_index; // @[SIMT_STACK.scala 160:{29,29}]
  wire  ipdom_index_1 = ~ipdom_stack_4_1_index; // @[SIMT_STACK.scala 229:28]
  wire  _push_2_T_3 = 2'h2 == warp_id; // @[SIMT_STACK.scala 200:75]
  wire  ipdom_stack_4_2_index = ipdom_stack_2_io_index; // @[SIMT_STACK.scala 160:{29,29}]
  wire  ipdom_index_2 = ~ipdom_stack_4_2_index; // @[SIMT_STACK.scala 229:28]
  wire  _push_3_T_3 = 2'h3 == warp_id; // @[SIMT_STACK.scala 200:75]
  wire  ipdom_stack_4_3_index = ipdom_stack_3_io_index; // @[SIMT_STACK.scala 160:{29,29}]
  wire  ipdom_index_3 = ~ipdom_stack_4_3_index; // @[SIMT_STACK.scala 229:28]
  wire [39:0] ipdom_stack_4_0_d = ipdom_stack_io_d; // @[SIMT_STACK.scala 160:{29,29}]
  wire [39:0] ipdom_stack_4_1_d = ipdom_stack_1_io_d; // @[SIMT_STACK.scala 160:{29,29}]
  wire [39:0] _GEN_10 = 2'h1 == warp_id ? ipdom_stack_4_1_d : ipdom_stack_4_0_d; // @[SIMT_STACK.scala 242:{36,36}]
  wire [39:0] ipdom_stack_4_2_d = ipdom_stack_2_io_d; // @[SIMT_STACK.scala 160:{29,29}]
  wire [39:0] _GEN_11 = 2'h2 == warp_id ? ipdom_stack_4_2_d : _GEN_10; // @[SIMT_STACK.scala 242:{36,36}]
  wire [39:0] ipdom_stack_4_3_d = ipdom_stack_3_io_d; // @[SIMT_STACK.scala 160:{29,29}]
  wire [39:0] _GEN_12 = 2'h3 == warp_id ? ipdom_stack_4_3_d : _GEN_11; // @[SIMT_STACK.scala 242:{36,36}]
  wire [31:0] join_pc = _GEN_12[39:8]; // @[SIMT_STACK.scala 242:36]
  wire [7:0] join_tm = _GEN_12[7:0]; // @[SIMT_STACK.scala 243:36]
  wire  _GEN_14 = 2'h1 == warp_id ? ipdom_index_1 : ipdom_index_0; // @[SIMT_STACK.scala 244:{13,13}]
  wire  _GEN_15 = 2'h2 == warp_id ? ipdom_index_2 : _GEN_14; // @[SIMT_STACK.scala 244:{13,13}]
  wire  join_index = 2'h3 == warp_id ? ipdom_index_3 : _GEN_15; // @[SIMT_STACK.scala 244:{13,13}]
  wire  ipdom_stack_4_0_pairo = ipdom_stack_io_pairo; // @[SIMT_STACK.scala 160:{29,29}]
  wire  ipdom_stack_4_1_pairo = ipdom_stack_1_io_pairo; // @[SIMT_STACK.scala 160:{29,29}]
  wire  _GEN_18 = 2'h1 == warp_id ? ipdom_stack_4_1_pairo : ipdom_stack_4_0_pairo; // @[SIMT_STACK.scala 245:{13,13}]
  wire  ipdom_stack_4_2_pairo = ipdom_stack_2_io_pairo; // @[SIMT_STACK.scala 160:{29,29}]
  wire  _GEN_19 = 2'h2 == warp_id ? ipdom_stack_4_2_pairo : _GEN_18; // @[SIMT_STACK.scala 245:{13,13}]
  wire  ipdom_stack_4_3_pairo = ipdom_stack_3_io_pairo; // @[SIMT_STACK.scala 160:{29,29}]
  wire  join_pair = 2'h3 == warp_id ? ipdom_stack_4_3_pairo : _GEN_19; // @[SIMT_STACK.scala 245:{13,13}]
  wire  _T_8 = opcode & branch_ctl_buf_io_deq_valid; // @[SIMT_STACK.scala 256:23]
  wire  _T_10 = ~join_pair; // @[SIMT_STACK.scala 260:16]
  wire [31:0] _GEN_22 = ~join_pair ? branch_ctl_buf_io_deq_bits_PC_branch : 32'h0; // @[SIMT_STACK.scala 253:20 260:27 262:24]
  wire [31:0] _GEN_23 = join_index ? join_pc : _GEN_22; // @[SIMT_STACK.scala 257:29 258:24]
  wire  _GEN_24 = join_index | _T_10; // @[SIMT_STACK.scala 257:29 259:22]
  wire  _GEN_26 = elseOnly & branch_ctl_buf_io_deq_valid; // @[SIMT_STACK.scala 255:19 267:19 269:23]
  wire [1:0] _GEN_27 = elseOnly ? warp_id : 2'h0; // @[SIMT_STACK.scala 252:17 267:19 270:21]
  wire [31:0] _GEN_28 = elseOnly ? branch_ctl_buf_io_deq_bits_PC_branch : 32'h0; // @[SIMT_STACK.scala 267:19 253:20 271:24]
  wire  _GEN_29 = _T & branch_ctl_buf_io_deq_valid & elseOnly; // @[SIMT_STACK.scala 254:18 266:53]
  wire  _GEN_30 = _T & branch_ctl_buf_io_deq_valid & _GEN_26; // @[SIMT_STACK.scala 255:19 266:53]
  wire [1:0] _GEN_31 = _T & branch_ctl_buf_io_deq_valid ? _GEN_27 : 2'h0; // @[SIMT_STACK.scala 252:17 266:53]
  wire [31:0] _GEN_32 = _T & branch_ctl_buf_io_deq_valid ? _GEN_28 : 32'h0; // @[SIMT_STACK.scala 253:20 266:53]
  wire [7:0] _GEN_62 = 2'h1 == io_input_wid ? thread_masks_1 : thread_masks_0; // @[SIMT_STACK.scala 289:{16,16}]
  wire [7:0] _GEN_63 = 2'h2 == io_input_wid ? thread_masks_2 : _GEN_62; // @[SIMT_STACK.scala 289:{16,16}]
  Queue_46 branch_ctl_buf ( // @[Decoupled.scala 361:21]
    .clock(branch_ctl_buf_clock),
    .reset(branch_ctl_buf_reset),
    .io_enq_ready(branch_ctl_buf_io_enq_ready),
    .io_enq_valid(branch_ctl_buf_io_enq_valid),
    .io_enq_bits_opcode(branch_ctl_buf_io_enq_bits_opcode),
    .io_enq_bits_wid(branch_ctl_buf_io_enq_bits_wid),
    .io_enq_bits_PC_branch(branch_ctl_buf_io_enq_bits_PC_branch),
    .io_enq_bits_mask_init(branch_ctl_buf_io_enq_bits_mask_init),
    .io_deq_ready(branch_ctl_buf_io_deq_ready),
    .io_deq_valid(branch_ctl_buf_io_deq_valid),
    .io_deq_bits_opcode(branch_ctl_buf_io_deq_bits_opcode),
    .io_deq_bits_wid(branch_ctl_buf_io_deq_bits_wid),
    .io_deq_bits_PC_branch(branch_ctl_buf_io_deq_bits_PC_branch),
    .io_deq_bits_mask_init(branch_ctl_buf_io_deq_bits_mask_init)
  );
  Queue_47 fetch_ctl_buf ( // @[SIMT_STACK.scala 133:29]
    .clock(fetch_ctl_buf_clock),
    .reset(fetch_ctl_buf_reset),
    .io_enq_ready(fetch_ctl_buf_io_enq_ready),
    .io_enq_valid(fetch_ctl_buf_io_enq_valid),
    .io_enq_bits_wid(fetch_ctl_buf_io_enq_bits_wid),
    .io_enq_bits_jump(fetch_ctl_buf_io_enq_bits_jump),
    .io_enq_bits_new_pc(fetch_ctl_buf_io_enq_bits_new_pc),
    .io_deq_ready(fetch_ctl_buf_io_deq_ready),
    .io_deq_valid(fetch_ctl_buf_io_deq_valid),
    .io_deq_bits_wid(fetch_ctl_buf_io_deq_bits_wid),
    .io_deq_bits_jump(fetch_ctl_buf_io_deq_bits_jump),
    .io_deq_bits_new_pc(fetch_ctl_buf_io_deq_bits_new_pc)
  );
  ipdom_stack ipdom_stack ( // @[SIMT_STACK.scala 160:55]
    .clock(ipdom_stack_clock),
    .reset(ipdom_stack_reset),
    .io_push(ipdom_stack_io_push),
    .io_pop(ipdom_stack_io_pop),
    .io_pair(ipdom_stack_io_pair),
    .io_branchImm(ipdom_stack_io_branchImm),
    .io_q1(ipdom_stack_io_q1),
    .io_q2(ipdom_stack_io_q2),
    .io_d(ipdom_stack_io_d),
    .io_index(ipdom_stack_io_index),
    .io_pairo(ipdom_stack_io_pairo)
  );
  ipdom_stack ipdom_stack_1 ( // @[SIMT_STACK.scala 160:55]
    .clock(ipdom_stack_1_clock),
    .reset(ipdom_stack_1_reset),
    .io_push(ipdom_stack_1_io_push),
    .io_pop(ipdom_stack_1_io_pop),
    .io_pair(ipdom_stack_1_io_pair),
    .io_branchImm(ipdom_stack_1_io_branchImm),
    .io_q1(ipdom_stack_1_io_q1),
    .io_q2(ipdom_stack_1_io_q2),
    .io_d(ipdom_stack_1_io_d),
    .io_index(ipdom_stack_1_io_index),
    .io_pairo(ipdom_stack_1_io_pairo)
  );
  ipdom_stack ipdom_stack_2 ( // @[SIMT_STACK.scala 160:55]
    .clock(ipdom_stack_2_clock),
    .reset(ipdom_stack_2_reset),
    .io_push(ipdom_stack_2_io_push),
    .io_pop(ipdom_stack_2_io_pop),
    .io_pair(ipdom_stack_2_io_pair),
    .io_branchImm(ipdom_stack_2_io_branchImm),
    .io_q1(ipdom_stack_2_io_q1),
    .io_q2(ipdom_stack_2_io_q2),
    .io_d(ipdom_stack_2_io_d),
    .io_index(ipdom_stack_2_io_index),
    .io_pairo(ipdom_stack_2_io_pairo)
  );
  ipdom_stack ipdom_stack_3 ( // @[SIMT_STACK.scala 160:55]
    .clock(ipdom_stack_3_clock),
    .reset(ipdom_stack_3_reset),
    .io_push(ipdom_stack_3_io_push),
    .io_pop(ipdom_stack_3_io_pop),
    .io_pair(ipdom_stack_3_io_pair),
    .io_branchImm(ipdom_stack_3_io_branchImm),
    .io_q1(ipdom_stack_3_io_q1),
    .io_q2(ipdom_stack_3_io_q2),
    .io_d(ipdom_stack_3_io_d),
    .io_index(ipdom_stack_3_io_index),
    .io_pairo(ipdom_stack_3_io_pairo)
  );
  assign io_branch_ctl_ready = branch_ctl_buf_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_if_mask_ready = fetch_ctl_buf_io_enq_ready; // @[Decoupled.scala 355:21 SIMT_STACK.scala 195:21]
  assign io_out_mask = 2'h3 == io_input_wid ? thread_masks_3 : _GEN_63; // @[SIMT_STACK.scala 289:{16,16}]
  assign io_complete_valid = _branch_ctl_buf_io_deq_ready_T & _T & branch_ctl_buf_io_deq_valid & ~elseOnly; // @[SIMT_STACK.scala 196:75]
  assign io_complete_bits = branch_ctl_buf_io_deq_bits_wid; // @[SIMT_STACK.scala 197:19]
  assign io_fetch_ctl_valid = fetch_ctl_buf_io_deq_valid; // @[SIMT_STACK.scala 277:16]
  assign io_fetch_ctl_bits_wid = fetch_ctl_buf_io_deq_bits_wid; // @[SIMT_STACK.scala 277:16]
  assign io_fetch_ctl_bits_jump = fetch_ctl_buf_io_deq_bits_jump; // @[SIMT_STACK.scala 277:16]
  assign io_fetch_ctl_bits_new_pc = fetch_ctl_buf_io_deq_bits_new_pc; // @[SIMT_STACK.scala 277:16]
  assign branch_ctl_buf_clock = clock;
  assign branch_ctl_buf_reset = reset;
  assign branch_ctl_buf_io_enq_valid = io_branch_ctl_valid; // @[Decoupled.scala 363:22]
  assign branch_ctl_buf_io_enq_bits_opcode = io_branch_ctl_bits_opcode; // @[Decoupled.scala 364:21]
  assign branch_ctl_buf_io_enq_bits_wid = io_branch_ctl_bits_wid; // @[Decoupled.scala 364:21]
  assign branch_ctl_buf_io_enq_bits_PC_branch = io_branch_ctl_bits_PC_branch; // @[Decoupled.scala 364:21]
  assign branch_ctl_buf_io_enq_bits_mask_init = io_branch_ctl_bits_mask_init; // @[Decoupled.scala 364:21]
  assign branch_ctl_buf_io_deq_ready = fetch_ctl_buf_io_enq_ready & _GEN_1; // @[SIMT_STACK.scala 165:35 182:26]
  assign fetch_ctl_buf_clock = clock;
  assign fetch_ctl_buf_reset = reset;
  assign fetch_ctl_buf_io_enq_valid = opcode & branch_ctl_buf_io_deq_valid ? branch_ctl_buf_io_deq_valid : _GEN_30; // @[SIMT_STACK.scala 256:47 264:21]
  assign fetch_ctl_buf_io_enq_bits_wid = opcode & branch_ctl_buf_io_deq_valid ? warp_id : _GEN_31; // @[SIMT_STACK.scala 256:47 265:19]
  assign fetch_ctl_buf_io_enq_bits_jump = opcode & branch_ctl_buf_io_deq_valid ? _GEN_24 : _GEN_29; // @[SIMT_STACK.scala 256:47]
  assign fetch_ctl_buf_io_enq_bits_new_pc = opcode & branch_ctl_buf_io_deq_valid ? _GEN_23 : _GEN_32; // @[SIMT_STACK.scala 256:47]
  assign fetch_ctl_buf_io_deq_ready = io_fetch_ctl_ready; // @[SIMT_STACK.scala 277:16]
  assign ipdom_stack_clock = clock;
  assign ipdom_stack_reset = reset;
  assign ipdom_stack_io_push = _T & _push_0_T_1 & 2'h0 == warp_id; // @[SIMT_STACK.scala 200:60]
  assign ipdom_stack_io_pop = opcode & _push_0_T_1 & _push_0_T_3; // @[SIMT_STACK.scala 201:60]
  assign ipdom_stack_io_pair = _branch_ctl_buf_io_deq_ready_T ? _diverge_T != 8'h0 : 1'h1; // @[SIMT_STACK.scala 188:12 190:28 192:13]
  assign ipdom_stack_io_branchImm = _branch_ctl_buf_io_deq_ready_T & else_mask == _GEN_6; // @[SIMT_STACK.scala 189:12 190:28 191:13]
  assign ipdom_stack_io_q1 = {32'h0,_GEN_6}; // @[Cat.scala 31:58]
  assign ipdom_stack_io_q2 = {PC_branch,_diverge_T}; // @[Cat.scala 31:58]
  assign ipdom_stack_1_clock = clock;
  assign ipdom_stack_1_reset = reset;
  assign ipdom_stack_1_io_push = _T & _push_0_T_1 & 2'h1 == warp_id; // @[SIMT_STACK.scala 200:60]
  assign ipdom_stack_1_io_pop = opcode & _push_0_T_1 & _push_1_T_3; // @[SIMT_STACK.scala 201:60]
  assign ipdom_stack_1_io_pair = _branch_ctl_buf_io_deq_ready_T ? _diverge_T != 8'h0 : 1'h1; // @[SIMT_STACK.scala 188:12 190:28 192:13]
  assign ipdom_stack_1_io_branchImm = _branch_ctl_buf_io_deq_ready_T & else_mask == _GEN_6; // @[SIMT_STACK.scala 189:12 190:28 191:13]
  assign ipdom_stack_1_io_q1 = {32'h0,_GEN_6}; // @[Cat.scala 31:58]
  assign ipdom_stack_1_io_q2 = {PC_branch,_diverge_T}; // @[Cat.scala 31:58]
  assign ipdom_stack_2_clock = clock;
  assign ipdom_stack_2_reset = reset;
  assign ipdom_stack_2_io_push = _T & _push_0_T_1 & 2'h2 == warp_id; // @[SIMT_STACK.scala 200:60]
  assign ipdom_stack_2_io_pop = opcode & _push_0_T_1 & _push_2_T_3; // @[SIMT_STACK.scala 201:60]
  assign ipdom_stack_2_io_pair = _branch_ctl_buf_io_deq_ready_T ? _diverge_T != 8'h0 : 1'h1; // @[SIMT_STACK.scala 188:12 190:28 192:13]
  assign ipdom_stack_2_io_branchImm = _branch_ctl_buf_io_deq_ready_T & else_mask == _GEN_6; // @[SIMT_STACK.scala 189:12 190:28 191:13]
  assign ipdom_stack_2_io_q1 = {32'h0,_GEN_6}; // @[Cat.scala 31:58]
  assign ipdom_stack_2_io_q2 = {PC_branch,_diverge_T}; // @[Cat.scala 31:58]
  assign ipdom_stack_3_clock = clock;
  assign ipdom_stack_3_reset = reset;
  assign ipdom_stack_3_io_push = _T & _push_0_T_1 & 2'h3 == warp_id; // @[SIMT_STACK.scala 200:60]
  assign ipdom_stack_3_io_pop = opcode & _push_0_T_1 & _push_3_T_3; // @[SIMT_STACK.scala 201:60]
  assign ipdom_stack_3_io_pair = _branch_ctl_buf_io_deq_ready_T ? _diverge_T != 8'h0 : 1'h1; // @[SIMT_STACK.scala 188:12 190:28 192:13]
  assign ipdom_stack_3_io_branchImm = _branch_ctl_buf_io_deq_ready_T & else_mask == _GEN_6; // @[SIMT_STACK.scala 189:12 190:28 191:13]
  assign ipdom_stack_3_io_q1 = {32'h0,_GEN_6}; // @[Cat.scala 31:58]
  assign ipdom_stack_3_io_q2 = {PC_branch,_diverge_T}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[SIMT_STACK.scala 137:29]
      thread_masks_0 <= 8'hff; // @[SIMT_STACK.scala 137:29]
    end else if (_branch_ctl_buf_io_deq_ready_T) begin // @[SIMT_STACK.scala 279:27]
      if (_io_complete_valid_T_4) begin // @[SIMT_STACK.scala 280:21]
        if (2'h0 == warp_id) begin // @[SIMT_STACK.scala 281:29]
          thread_masks_0 <= if_mask; // @[SIMT_STACK.scala 281:29]
        end
      end else if (2'h0 == warp_id) begin // @[SIMT_STACK.scala 283:29]
        thread_masks_0 <= _diverge_T; // @[SIMT_STACK.scala 283:29]
      end
    end else if (_T_8) begin // @[SIMT_STACK.scala 285:52]
      if (2'h0 == warp_id) begin // @[SIMT_STACK.scala 286:27]
        thread_masks_0 <= join_tm; // @[SIMT_STACK.scala 286:27]
      end
    end
    if (reset) begin // @[SIMT_STACK.scala 137:29]
      thread_masks_1 <= 8'hff; // @[SIMT_STACK.scala 137:29]
    end else if (_branch_ctl_buf_io_deq_ready_T) begin // @[SIMT_STACK.scala 279:27]
      if (_io_complete_valid_T_4) begin // @[SIMT_STACK.scala 280:21]
        if (2'h1 == warp_id) begin // @[SIMT_STACK.scala 281:29]
          thread_masks_1 <= if_mask; // @[SIMT_STACK.scala 281:29]
        end
      end else if (2'h1 == warp_id) begin // @[SIMT_STACK.scala 283:29]
        thread_masks_1 <= _diverge_T; // @[SIMT_STACK.scala 283:29]
      end
    end else if (_T_8) begin // @[SIMT_STACK.scala 285:52]
      if (2'h1 == warp_id) begin // @[SIMT_STACK.scala 286:27]
        thread_masks_1 <= join_tm; // @[SIMT_STACK.scala 286:27]
      end
    end
    if (reset) begin // @[SIMT_STACK.scala 137:29]
      thread_masks_2 <= 8'hff; // @[SIMT_STACK.scala 137:29]
    end else if (_branch_ctl_buf_io_deq_ready_T) begin // @[SIMT_STACK.scala 279:27]
      if (_io_complete_valid_T_4) begin // @[SIMT_STACK.scala 280:21]
        if (2'h2 == warp_id) begin // @[SIMT_STACK.scala 281:29]
          thread_masks_2 <= if_mask; // @[SIMT_STACK.scala 281:29]
        end
      end else if (2'h2 == warp_id) begin // @[SIMT_STACK.scala 283:29]
        thread_masks_2 <= _diverge_T; // @[SIMT_STACK.scala 283:29]
      end
    end else if (_T_8) begin // @[SIMT_STACK.scala 285:52]
      if (2'h2 == warp_id) begin // @[SIMT_STACK.scala 286:27]
        thread_masks_2 <= join_tm; // @[SIMT_STACK.scala 286:27]
      end
    end
    if (reset) begin // @[SIMT_STACK.scala 137:29]
      thread_masks_3 <= 8'hff; // @[SIMT_STACK.scala 137:29]
    end else if (_branch_ctl_buf_io_deq_ready_T) begin // @[SIMT_STACK.scala 279:27]
      if (_io_complete_valid_T_4) begin // @[SIMT_STACK.scala 280:21]
        if (2'h3 == warp_id) begin // @[SIMT_STACK.scala 281:29]
          thread_masks_3 <= if_mask; // @[SIMT_STACK.scala 281:29]
        end
      end else if (2'h3 == warp_id) begin // @[SIMT_STACK.scala 283:29]
        thread_masks_3 <= _diverge_T; // @[SIMT_STACK.scala 283:29]
      end
    end else if (_T_8) begin // @[SIMT_STACK.scala 285:52]
      if (2'h3 == warp_id) begin // @[SIMT_STACK.scala 286:27]
        thread_masks_3 <= join_tm; // @[SIMT_STACK.scala 286:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  thread_masks_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  thread_masks_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  thread_masks_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  thread_masks_3 = _RAND_3[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_13(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_wid,
  input         io_in_0_bits_jump,
  input  [31:0] io_in_0_bits_new_pc,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_wid,
  input         io_in_1_bits_jump,
  input  [31:0] io_in_1_bits_new_pc,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_wid,
  output        io_out_bits_jump,
  output [31:0] io_out_bits_new_pc
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_wid = io_in_0_valid ? io_in_0_bits_wid : io_in_1_bits_wid; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_jump = io_in_0_valid ? io_in_0_bits_jump : io_in_1_bits_jump; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_new_pc = io_in_0_valid ? io_in_0_bits_new_pc : io_in_1_bits_new_pc; // @[Arbiter.scala 139:15 141:26 143:19]
endmodule
module Branch_back(
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_wid,
  output        io_out_bits_jump,
  output [31:0] io_out_bits_new_pc,
  output        io_in0_ready,
  input         io_in0_valid,
  input  [1:0]  io_in0_bits_wid,
  input         io_in0_bits_jump,
  input  [31:0] io_in0_bits_new_pc,
  output        io_in1_ready,
  input         io_in1_valid,
  input  [1:0]  io_in1_bits_wid,
  input         io_in1_bits_jump,
  input  [31:0] io_in1_bits_new_pc
);
  wire  arbiter_io_in_0_ready; // @[writeback.scala 13:21]
  wire  arbiter_io_in_0_valid; // @[writeback.scala 13:21]
  wire [1:0] arbiter_io_in_0_bits_wid; // @[writeback.scala 13:21]
  wire  arbiter_io_in_0_bits_jump; // @[writeback.scala 13:21]
  wire [31:0] arbiter_io_in_0_bits_new_pc; // @[writeback.scala 13:21]
  wire  arbiter_io_in_1_ready; // @[writeback.scala 13:21]
  wire  arbiter_io_in_1_valid; // @[writeback.scala 13:21]
  wire [1:0] arbiter_io_in_1_bits_wid; // @[writeback.scala 13:21]
  wire  arbiter_io_in_1_bits_jump; // @[writeback.scala 13:21]
  wire [31:0] arbiter_io_in_1_bits_new_pc; // @[writeback.scala 13:21]
  wire  arbiter_io_out_ready; // @[writeback.scala 13:21]
  wire  arbiter_io_out_valid; // @[writeback.scala 13:21]
  wire [1:0] arbiter_io_out_bits_wid; // @[writeback.scala 13:21]
  wire  arbiter_io_out_bits_jump; // @[writeback.scala 13:21]
  wire [31:0] arbiter_io_out_bits_new_pc; // @[writeback.scala 13:21]
  Arbiter_13 arbiter ( // @[writeback.scala 13:21]
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_wid(arbiter_io_in_0_bits_wid),
    .io_in_0_bits_jump(arbiter_io_in_0_bits_jump),
    .io_in_0_bits_new_pc(arbiter_io_in_0_bits_new_pc),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_wid(arbiter_io_in_1_bits_wid),
    .io_in_1_bits_jump(arbiter_io_in_1_bits_jump),
    .io_in_1_bits_new_pc(arbiter_io_in_1_bits_new_pc),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_wid(arbiter_io_out_bits_wid),
    .io_out_bits_jump(arbiter_io_out_bits_jump),
    .io_out_bits_new_pc(arbiter_io_out_bits_new_pc)
  );
  assign io_out_valid = arbiter_io_out_valid; // @[writeback.scala 16:17]
  assign io_out_bits_wid = arbiter_io_out_bits_wid; // @[writeback.scala 16:17]
  assign io_out_bits_jump = arbiter_io_out_bits_jump; // @[writeback.scala 16:17]
  assign io_out_bits_new_pc = arbiter_io_out_bits_new_pc; // @[writeback.scala 16:17]
  assign io_in0_ready = arbiter_io_in_0_ready; // @[Decoupled.scala 355:21 writeback.scala 14:19]
  assign io_in1_ready = arbiter_io_in_1_ready; // @[Decoupled.scala 355:21 writeback.scala 15:19]
  assign arbiter_io_in_0_valid = io_in0_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_io_in_0_bits_wid = io_in0_bits_wid; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_io_in_0_bits_jump = io_in0_bits_jump; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_io_in_0_bits_new_pc = io_in0_bits_new_pc; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_io_in_1_valid = io_in1_valid; // @[Decoupled.scala 355:21 356:17]
  assign arbiter_io_in_1_bits_wid = io_in1_bits_wid; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_io_in_1_bits_jump = io_in1_bits_jump; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_io_in_1_bits_new_pc = io_in1_bits_new_pc; // @[Decoupled.scala 355:21 357:16]
  assign arbiter_io_out_ready = io_out_ready; // @[writeback.scala 16:17]
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input  [31:0] io_ctrl_inst,
  input  [1:0]  io_ctrl_csr,
  input         io_ctrl_isvec,
  input  [31:0] io_in1,
  input         io_write,
  output [31:0] io_wb_wxd_rd,
  output [2:0]  io_frm,
  input         io_CTA2csr_valid,
  input  [2:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count,
  input  [9:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch,
  input  [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch,
  input  [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch,
  input  [4:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch,
  input  [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  reg  MTIP; // @[CSR.scala 86:21]
  reg  MTIE; // @[CSR.scala 89:21]
  reg  MSIP; // @[CSR.scala 92:21]
  reg  MSIE; // @[CSR.scala 95:21]
  reg  MEIP; // @[CSR.scala 98:21]
  reg  MEIE; // @[CSR.scala 101:21]
  wire [31:0] mip = {20'h0,MEIP,2'h0,1'h0,MTIP,1'h0,2'h0,MSIP,3'h0}; // @[Cat.scala 31:58]
  wire [31:0] mie = {20'h0,MEIE,2'h0,1'h0,MTIE,1'h0,2'h0,MSIE,3'h0}; // @[Cat.scala 31:58]
  reg  MIE; // @[CSR.scala 107:21]
  reg  MPIE; // @[CSR.scala 110:21]
  wire [31:0] mstatus = {21'h3,3'h0,MPIE,2'h0,1'h0,MIE,1'h0,2'h0}; // @[Cat.scala 31:58]
  reg [31:0] mscratch; // @[CSR.scala 127:25]
  reg [31:0] mepc; // @[CSR.scala 130:21]
  reg [31:0] mcause; // @[CSR.scala 133:23]
  reg [31:0] mtval; // @[CSR.scala 136:22]
  reg [31:0] threadid; // @[CSR.scala 139:25]
  reg [2:0] wg_wf_count; // @[CSR.scala 143:24]
  reg [9:0] wf_size_dispatch; // @[CSR.scala 144:29]
  reg [12:0] sgpr_base_dispatch; // @[CSR.scala 145:31]
  reg [12:0] vgpr_base_dispatch; // @[CSR.scala 146:31]
  reg [4:0] wf_tag_dispatch; // @[CSR.scala 147:28]
  reg [12:0] lds_base_dispatch; // @[CSR.scala 148:30]
  reg  NV; // @[CSR.scala 152:19]
  reg  DZ; // @[CSR.scala 153:19]
  reg  OF; // @[CSR.scala 154:19]
  reg  UF; // @[CSR.scala 155:19]
  reg  NX; // @[CSR.scala 156:19]
  wire [4:0] fflags = {NV,DZ,OF,UF,NX}; // @[Cat.scala 31:58]
  reg [2:0] frm; // @[CSR.scala 158:20]
  wire [31:0] fcsr = {24'h0,frm,NV,DZ,OF,UF,NX}; // @[Cat.scala 31:58]
  wire [11:0] csr_addr = io_ctrl_inst[31:20]; // @[CSR.scala 177:30]
  wire  wen = |io_ctrl_csr & io_write; // @[CSR.scala 185:28]
  wire  _csr_rdata_T_1 = 12'h300 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_3 = 12'h304 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_5 = 12'h305 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_7 = 12'h340 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_9 = 12'h341 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_11 = 12'h342 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_13 = 12'h343 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_15 = 12'h344 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_17 = 12'h2 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_19 = 12'h3 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_21 = 12'h1 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_23 = 12'h800 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_25 = 12'hc21 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_27 = 12'h801 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_29 = 12'h802 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_31 = 12'h803 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_33 = 12'h804 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_35 = 12'h805 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_37 = 12'h806 == csr_addr; // @[Lookup.scala 31:38]
  wire  _csr_rdata_T_39 = 12'h807 == csr_addr; // @[Lookup.scala 31:38]
  wire [31:0] _csr_rdata_T_40 = _csr_rdata_T_39 ? 32'h1000 : 32'h0; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_41 = _csr_rdata_T_37 ? {{19'd0}, lds_base_dispatch} : _csr_rdata_T_40; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_42 = _csr_rdata_T_35 ? {{27'd0}, wf_tag_dispatch} : _csr_rdata_T_41; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_43 = _csr_rdata_T_33 ? {{19'd0}, vgpr_base_dispatch} : _csr_rdata_T_42; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_44 = _csr_rdata_T_31 ? {{19'd0}, sgpr_base_dispatch} : _csr_rdata_T_43; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_45 = _csr_rdata_T_29 ? {{22'd0}, wf_size_dispatch} : _csr_rdata_T_44; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_46 = _csr_rdata_T_27 ? {{29'd0}, wg_wf_count} : _csr_rdata_T_45; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_47 = _csr_rdata_T_25 ? 32'h10 : _csr_rdata_T_46; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_48 = _csr_rdata_T_23 ? threadid : _csr_rdata_T_47; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_49 = _csr_rdata_T_21 ? {{27'd0}, fflags} : _csr_rdata_T_48; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_50 = _csr_rdata_T_19 ? fcsr : _csr_rdata_T_49; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_51 = _csr_rdata_T_17 ? {{29'd0}, frm} : _csr_rdata_T_50; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_52 = _csr_rdata_T_15 ? mip : _csr_rdata_T_51; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_53 = _csr_rdata_T_13 ? mtval : _csr_rdata_T_52; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_54 = _csr_rdata_T_11 ? mcause : _csr_rdata_T_53; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_55 = _csr_rdata_T_9 ? mepc : _csr_rdata_T_54; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_56 = _csr_rdata_T_7 ? mscratch : _csr_rdata_T_55; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_57 = _csr_rdata_T_5 ? 32'h0 : _csr_rdata_T_56; // @[Lookup.scala 34:39]
  wire [31:0] _csr_rdata_T_58 = _csr_rdata_T_3 ? mie : _csr_rdata_T_57; // @[Lookup.scala 34:39]
  wire [31:0] csr_rdata = _csr_rdata_T_1 ? mstatus : _csr_rdata_T_58; // @[Lookup.scala 34:39]
  wire [31:0] _csr_wdata_T = csr_rdata | io_in1; // @[CSR.scala 186:92]
  wire [31:0] _csr_wdata_T_1 = ~io_in1; // @[CSR.scala 186:130]
  wire [31:0] _csr_wdata_T_2 = csr_rdata & _csr_wdata_T_1; // @[CSR.scala 186:127]
  wire [31:0] _csr_wdata_T_4 = 2'h1 == io_ctrl_csr ? io_in1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _csr_wdata_T_6 = 2'h2 == io_ctrl_csr ? _csr_wdata_T : _csr_wdata_T_4; // @[Mux.scala 81:58]
  wire [31:0] csr_wdata = 2'h3 == io_ctrl_csr ? _csr_wdata_T_2 : _csr_wdata_T_6; // @[Mux.scala 81:58]
  wire [32:0] _GEN_115 = {{1'd0}, io_in1}; // @[CSR.scala 218:23]
  wire [31:0] _wdata_T_3 = {{1'd0}, io_in1[31:1]}; // @[CSR.scala 218:55]
  wire [31:0] _wdata_T_4 = _GEN_115 > 33'h10 ? 32'h8 : _wdata_T_3; // @[CSR.scala 218:19]
  wire [31:0] _wdata_T_5 = io_in1 < 32'h8 ? io_in1 : _wdata_T_4; // @[CSR.scala 217:19]
  wire [31:0] _GEN_0 = csr_addr == 12'h343 ? csr_wdata : mtval; // @[CSR.scala 244:43 245:15 136:22]
  wire [31:0] _GEN_1 = csr_addr == 12'h342 ? csr_wdata : mcause; // @[CSR.scala 242:44 243:16 133:23]
  wire [31:0] _GEN_2 = csr_addr == 12'h342 ? mtval : _GEN_0; // @[CSR.scala 136:22 242:44]
  wire [31:0] _GEN_3 = csr_addr == 12'h341 ? csr_wdata : mepc; // @[CSR.scala 240:42 241:14 130:21]
  wire [31:0] _GEN_4 = csr_addr == 12'h341 ? mcause : _GEN_1; // @[CSR.scala 133:23 240:42]
  wire [31:0] _GEN_5 = csr_addr == 12'h341 ? mtval : _GEN_2; // @[CSR.scala 136:22 240:42]
  wire [31:0] _GEN_6 = csr_addr == 12'h340 ? csr_wdata : mscratch; // @[CSR.scala 238:46 239:18 127:25]
  wire [31:0] _GEN_7 = csr_addr == 12'h340 ? mepc : _GEN_3; // @[CSR.scala 130:21 238:46]
  wire [31:0] _GEN_8 = csr_addr == 12'h340 ? mcause : _GEN_4; // @[CSR.scala 133:23 238:46]
  wire [31:0] _GEN_9 = csr_addr == 12'h340 ? mtval : _GEN_5; // @[CSR.scala 136:22 238:46]
  wire  _GEN_10 = csr_addr == 12'h304 ? csr_wdata[7] : MTIE; // @[CSR.scala 234:42 235:14 89:21]
  wire  _GEN_11 = csr_addr == 12'h304 ? csr_wdata[3] : MSIE; // @[CSR.scala 234:42 236:14 95:21]
  wire  _GEN_12 = csr_addr == 12'h304 ? csr_wdata[11] : MEIE; // @[CSR.scala 234:42 237:14 101:21]
  wire [31:0] _GEN_13 = csr_addr == 12'h304 ? mscratch : _GEN_6; // @[CSR.scala 127:25 234:42]
  wire [31:0] _GEN_14 = csr_addr == 12'h304 ? mepc : _GEN_7; // @[CSR.scala 130:21 234:42]
  wire [31:0] _GEN_15 = csr_addr == 12'h304 ? mcause : _GEN_8; // @[CSR.scala 133:23 234:42]
  wire [31:0] _GEN_16 = csr_addr == 12'h304 ? mtval : _GEN_9; // @[CSR.scala 136:22 234:42]
  wire  _GEN_17 = csr_addr == 12'h344 ? csr_wdata[7] : MTIP; // @[CSR.scala 230:42 231:14 86:21]
  wire  _GEN_18 = csr_addr == 12'h344 ? csr_wdata[3] : MSIP; // @[CSR.scala 230:42 232:14 92:21]
  wire  _GEN_19 = csr_addr == 12'h344 ? csr_wdata[11] : MEIP; // @[CSR.scala 230:42 233:14 98:21]
  wire  _GEN_20 = csr_addr == 12'h344 ? MTIE : _GEN_10; // @[CSR.scala 230:42 89:21]
  wire  _GEN_21 = csr_addr == 12'h344 ? MSIE : _GEN_11; // @[CSR.scala 230:42 95:21]
  wire  _GEN_22 = csr_addr == 12'h344 ? MEIE : _GEN_12; // @[CSR.scala 101:21 230:42]
  wire [31:0] _GEN_23 = csr_addr == 12'h344 ? mscratch : _GEN_13; // @[CSR.scala 127:25 230:42]
  wire [31:0] _GEN_24 = csr_addr == 12'h344 ? mepc : _GEN_14; // @[CSR.scala 130:21 230:42]
  wire [31:0] _GEN_25 = csr_addr == 12'h344 ? mcause : _GEN_15; // @[CSR.scala 133:23 230:42]
  wire [31:0] _GEN_26 = csr_addr == 12'h344 ? mtval : _GEN_16; // @[CSR.scala 136:22 230:42]
  wire  _GEN_27 = csr_addr == 12'h300 ? csr_wdata[3] : MIE; // @[CSR.scala 227:46 228:13 107:21]
  wire  _GEN_28 = csr_addr == 12'h300 ? csr_wdata[7] : MPIE; // @[CSR.scala 227:46 229:14 110:21]
  wire  _GEN_29 = csr_addr == 12'h300 ? MTIP : _GEN_17; // @[CSR.scala 227:46 86:21]
  wire  _GEN_30 = csr_addr == 12'h300 ? MSIP : _GEN_18; // @[CSR.scala 227:46 92:21]
  wire  _GEN_31 = csr_addr == 12'h300 ? MEIP : _GEN_19; // @[CSR.scala 227:46 98:21]
  wire  _GEN_32 = csr_addr == 12'h300 ? MTIE : _GEN_20; // @[CSR.scala 227:46 89:21]
  wire  _GEN_33 = csr_addr == 12'h300 ? MSIE : _GEN_21; // @[CSR.scala 227:46 95:21]
  wire  _GEN_34 = csr_addr == 12'h300 ? MEIE : _GEN_22; // @[CSR.scala 101:21 227:46]
  wire [31:0] _GEN_35 = csr_addr == 12'h300 ? mscratch : _GEN_23; // @[CSR.scala 127:25 227:46]
  wire [31:0] _GEN_36 = csr_addr == 12'h300 ? mepc : _GEN_24; // @[CSR.scala 130:21 227:46]
  wire [31:0] _GEN_37 = csr_addr == 12'h300 ? mcause : _GEN_25; // @[CSR.scala 133:23 227:46]
  wire [31:0] _GEN_38 = csr_addr == 12'h300 ? mtval : _GEN_26; // @[CSR.scala 136:22 227:46]
  wire [2:0] _GEN_39 = csr_addr == 12'h2 ? csr_wdata[2:0] : frm; // @[CSR.scala 225:41 226:12 158:20]
  wire  _GEN_40 = csr_addr == 12'h2 ? MIE : _GEN_27; // @[CSR.scala 107:21 225:41]
  wire  _GEN_41 = csr_addr == 12'h2 ? MPIE : _GEN_28; // @[CSR.scala 110:21 225:41]
  wire  _GEN_42 = csr_addr == 12'h2 ? MTIP : _GEN_29; // @[CSR.scala 225:41 86:21]
  wire  _GEN_43 = csr_addr == 12'h2 ? MSIP : _GEN_30; // @[CSR.scala 225:41 92:21]
  wire  _GEN_44 = csr_addr == 12'h2 ? MEIP : _GEN_31; // @[CSR.scala 225:41 98:21]
  wire  _GEN_45 = csr_addr == 12'h2 ? MTIE : _GEN_32; // @[CSR.scala 225:41 89:21]
  wire  _GEN_46 = csr_addr == 12'h2 ? MSIE : _GEN_33; // @[CSR.scala 225:41 95:21]
  wire  _GEN_47 = csr_addr == 12'h2 ? MEIE : _GEN_34; // @[CSR.scala 101:21 225:41]
  wire [31:0] _GEN_48 = csr_addr == 12'h2 ? mscratch : _GEN_35; // @[CSR.scala 127:25 225:41]
  wire [31:0] _GEN_49 = csr_addr == 12'h2 ? mepc : _GEN_36; // @[CSR.scala 130:21 225:41]
  wire [31:0] _GEN_50 = csr_addr == 12'h2 ? mcause : _GEN_37; // @[CSR.scala 133:23 225:41]
  wire [31:0] _GEN_51 = csr_addr == 12'h2 ? mtval : _GEN_38; // @[CSR.scala 136:22 225:41]
  wire [31:0] _GEN_70 = io_ctrl_isvec ? _wdata_T_5 : csr_rdata; // @[CSR.scala 216:26 217:14 182:8]
  wire [5:0] _threadid_T_1 = {io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch[2:0], 3'h0}; // @[CSR.scala 257:84]
  assign io_wb_wxd_rd = wen ? _GEN_70 : csr_rdata; // @[CSR.scala 215:14 182:8]
  assign io_frm = frm; // @[CSR.scala 160:9]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 86:21]
      MTIP <= 1'h0; // @[CSR.scala 86:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MTIP <= _GEN_42;
        end
      end
    end
    if (reset) begin // @[CSR.scala 89:21]
      MTIE <= 1'h0; // @[CSR.scala 89:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MTIE <= _GEN_45;
        end
      end
    end
    if (reset) begin // @[CSR.scala 92:21]
      MSIP <= 1'h0; // @[CSR.scala 92:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MSIP <= _GEN_43;
        end
      end
    end
    if (reset) begin // @[CSR.scala 95:21]
      MSIE <= 1'h0; // @[CSR.scala 95:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MSIE <= _GEN_46;
        end
      end
    end
    if (reset) begin // @[CSR.scala 98:21]
      MEIP <= 1'h0; // @[CSR.scala 98:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MEIP <= _GEN_44;
        end
      end
    end
    if (reset) begin // @[CSR.scala 101:21]
      MEIE <= 1'h0; // @[CSR.scala 101:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MEIE <= _GEN_47;
        end
      end
    end
    if (reset) begin // @[CSR.scala 107:21]
      MIE <= 1'h0; // @[CSR.scala 107:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MIE <= _GEN_40;
        end
      end
    end
    if (reset) begin // @[CSR.scala 110:21]
      MPIE <= 1'h0; // @[CSR.scala 110:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          MPIE <= _GEN_41;
        end
      end
    end
    if (reset) begin // @[CSR.scala 127:25]
      mscratch <= 32'h0; // @[CSR.scala 127:25]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          mscratch <= _GEN_48;
        end
      end
    end
    if (reset) begin // @[CSR.scala 130:21]
      mepc <= 32'h0; // @[CSR.scala 130:21]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          mepc <= _GEN_49;
        end
      end
    end
    if (reset) begin // @[CSR.scala 133:23]
      mcause <= 32'h0; // @[CSR.scala 133:23]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          mcause <= _GEN_50;
        end
      end
    end
    if (reset) begin // @[CSR.scala 136:22]
      mtval <= 32'h0; // @[CSR.scala 136:22]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          mtval <= _GEN_51;
        end
      end
    end
    if (reset) begin // @[CSR.scala 139:25]
      threadid <= 32'h0; // @[CSR.scala 139:25]
    end else if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      threadid <= {{26'd0}, _threadid_T_1}; // @[CSR.scala 257:13]
    end
    if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      wg_wf_count <= io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 250:17]
    end
    if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      wf_size_dispatch <= io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 251:22]
    end
    if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      sgpr_base_dispatch <= io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 252:23]
    end
    if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      vgpr_base_dispatch <= io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 253:23]
    end
    if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      wf_tag_dispatch <= io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 254:21]
    end
    if (io_CTA2csr_valid) begin // @[CSR.scala 248:25]
      lds_base_dispatch <= io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 255:22]
    end
    if (reset) begin // @[CSR.scala 152:19]
      NV <= 1'h0; // @[CSR.scala 152:19]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (csr_addr == 12'h1) begin // @[CSR.scala 219:43]
          NV <= csr_wdata[4]; // @[CSR.scala 224:11]
        end
      end
    end
    if (reset) begin // @[CSR.scala 153:19]
      DZ <= 1'h0; // @[CSR.scala 153:19]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (csr_addr == 12'h1) begin // @[CSR.scala 219:43]
          DZ <= csr_wdata[3]; // @[CSR.scala 223:11]
        end
      end
    end
    if (reset) begin // @[CSR.scala 154:19]
      OF <= 1'h0; // @[CSR.scala 154:19]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (csr_addr == 12'h1) begin // @[CSR.scala 219:43]
          OF <= csr_wdata[2]; // @[CSR.scala 222:11]
        end
      end
    end
    if (reset) begin // @[CSR.scala 155:19]
      UF <= 1'h0; // @[CSR.scala 155:19]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (csr_addr == 12'h1) begin // @[CSR.scala 219:43]
          UF <= csr_wdata[1]; // @[CSR.scala 221:11]
        end
      end
    end
    if (reset) begin // @[CSR.scala 156:19]
      NX <= 1'h0; // @[CSR.scala 156:19]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (csr_addr == 12'h1) begin // @[CSR.scala 219:43]
          NX <= csr_wdata[0]; // @[CSR.scala 220:11]
        end
      end
    end
    if (reset) begin // @[CSR.scala 158:20]
      frm <= 3'h0; // @[CSR.scala 158:20]
    end else if (wen) begin // @[CSR.scala 215:14]
      if (!(io_ctrl_isvec)) begin // @[CSR.scala 216:26]
        if (!(csr_addr == 12'h1)) begin // @[CSR.scala 219:43]
          frm <= _GEN_39;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  MTIP = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  MTIE = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  MSIP = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  MSIE = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  MEIP = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  MEIE = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  MIE = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  MPIE = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mscratch = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mepc = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mcause = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mtval = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  threadid = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  wg_wf_count = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  wf_size_dispatch = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  sgpr_base_dispatch = _RAND_15[12:0];
  _RAND_16 = {1{`RANDOM}};
  vgpr_base_dispatch = _RAND_16[12:0];
  _RAND_17 = {1{`RANDOM}};
  wf_tag_dispatch = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  lds_base_dispatch = _RAND_18[12:0];
  _RAND_19 = {1{`RANDOM}};
  NV = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  DZ = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  OF = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  UF = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  NX = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  frm = _RAND_24[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSRexe(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_ctrl_inst,
  input  [1:0]  io_in_bits_ctrl_wid,
  input  [1:0]  io_in_bits_ctrl_csr,
  input         io_in_bits_ctrl_isvec,
  input  [4:0]  io_in_bits_ctrl_reg_idxw,
  input         io_in_bits_ctrl_wxd,
  input  [31:0] io_in_bits_in1,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_wb_wxd_rd,
  output        io_out_bits_wxd,
  output [4:0]  io_out_bits_reg_idxw,
  output [1:0]  io_out_bits_warp_id,
  input  [1:0]  io_frm_wid,
  output [2:0]  io_frm,
  input         io_CTA2csr_valid,
  input  [2:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count,
  input  [9:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch,
  input  [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch,
  input  [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch,
  input  [4:0]  io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch,
  input  [12:0] io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch,
  input  [1:0]  io_CTA2csr_bits_wid
);
  wire  CSRFile_clock; // @[CSR.scala 270:45]
  wire  CSRFile_reset; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_io_ctrl_inst; // @[CSR.scala 270:45]
  wire [1:0] CSRFile_io_ctrl_csr; // @[CSR.scala 270:45]
  wire  CSRFile_io_ctrl_isvec; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_io_in1; // @[CSR.scala 270:45]
  wire  CSRFile_io_write; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_io_wb_wxd_rd; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_io_frm; // @[CSR.scala 270:45]
  wire  CSRFile_io_CTA2csr_valid; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:45]
  wire [9:0] CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [4:0] CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:45]
  wire  CSRFile_1_clock; // @[CSR.scala 270:45]
  wire  CSRFile_1_reset; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_1_io_ctrl_inst; // @[CSR.scala 270:45]
  wire [1:0] CSRFile_1_io_ctrl_csr; // @[CSR.scala 270:45]
  wire  CSRFile_1_io_ctrl_isvec; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_1_io_in1; // @[CSR.scala 270:45]
  wire  CSRFile_1_io_write; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_1_io_wb_wxd_rd; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_1_io_frm; // @[CSR.scala 270:45]
  wire  CSRFile_1_io_CTA2csr_valid; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:45]
  wire [9:0] CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [4:0] CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:45]
  wire  CSRFile_2_clock; // @[CSR.scala 270:45]
  wire  CSRFile_2_reset; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_2_io_ctrl_inst; // @[CSR.scala 270:45]
  wire [1:0] CSRFile_2_io_ctrl_csr; // @[CSR.scala 270:45]
  wire  CSRFile_2_io_ctrl_isvec; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_2_io_in1; // @[CSR.scala 270:45]
  wire  CSRFile_2_io_write; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_2_io_wb_wxd_rd; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_2_io_frm; // @[CSR.scala 270:45]
  wire  CSRFile_2_io_CTA2csr_valid; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:45]
  wire [9:0] CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [4:0] CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:45]
  wire  CSRFile_3_clock; // @[CSR.scala 270:45]
  wire  CSRFile_3_reset; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_3_io_ctrl_inst; // @[CSR.scala 270:45]
  wire [1:0] CSRFile_3_io_ctrl_csr; // @[CSR.scala 270:45]
  wire  CSRFile_3_io_ctrl_isvec; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_3_io_in1; // @[CSR.scala 270:45]
  wire  CSRFile_3_io_write; // @[CSR.scala 270:45]
  wire [31:0] CSRFile_3_io_wb_wxd_rd; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_3_io_frm; // @[CSR.scala 270:45]
  wire  CSRFile_3_io_CTA2csr_valid; // @[CSR.scala 270:45]
  wire [2:0] CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:45]
  wire [9:0] CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:45]
  wire [4:0] CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:45]
  wire [12:0] CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:45]
  wire  result_clock; // @[CSR.scala 280:20]
  wire  result_reset; // @[CSR.scala 280:20]
  wire  result_io_enq_ready; // @[CSR.scala 280:20]
  wire  result_io_enq_valid; // @[CSR.scala 280:20]
  wire [31:0] result_io_enq_bits_wb_wxd_rd; // @[CSR.scala 280:20]
  wire  result_io_enq_bits_wxd; // @[CSR.scala 280:20]
  wire [4:0] result_io_enq_bits_reg_idxw; // @[CSR.scala 280:20]
  wire [1:0] result_io_enq_bits_warp_id; // @[CSR.scala 280:20]
  wire  result_io_deq_ready; // @[CSR.scala 280:20]
  wire  result_io_deq_valid; // @[CSR.scala 280:20]
  wire [31:0] result_io_deq_bits_wb_wxd_rd; // @[CSR.scala 280:20]
  wire  result_io_deq_bits_wxd; // @[CSR.scala 280:20]
  wire [4:0] result_io_deq_bits_reg_idxw; // @[CSR.scala 280:20]
  wire [1:0] result_io_deq_bits_warp_id; // @[CSR.scala 280:20]
  wire  _vCSR_write_T = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  wire [31:0] vCSR_0_wb_wxd_rd = CSRFile_io_wb_wxd_rd; // @[CSR.scala 270:{19,19}]
  wire [31:0] vCSR_1_wb_wxd_rd = CSRFile_1_io_wb_wxd_rd; // @[CSR.scala 270:{19,19}]
  wire [31:0] _GEN_9 = 2'h1 == io_in_bits_ctrl_wid ? vCSR_1_wb_wxd_rd : vCSR_0_wb_wxd_rd; // @[CSR.scala 288:{31,31}]
  wire [31:0] vCSR_2_wb_wxd_rd = CSRFile_2_io_wb_wxd_rd; // @[CSR.scala 270:{19,19}]
  wire [31:0] _GEN_10 = 2'h2 == io_in_bits_ctrl_wid ? vCSR_2_wb_wxd_rd : _GEN_9; // @[CSR.scala 288:{31,31}]
  wire [31:0] vCSR_3_wb_wxd_rd = CSRFile_3_io_wb_wxd_rd; // @[CSR.scala 270:{19,19}]
  wire [2:0] vCSR_0_frm = CSRFile_io_frm; // @[CSR.scala 270:{19,19}]
  wire [2:0] vCSR_1_frm = CSRFile_1_io_frm; // @[CSR.scala 270:{19,19}]
  wire [2:0] _GEN_13 = 2'h1 == io_frm_wid ? vCSR_1_frm : vCSR_0_frm; // @[CSR.scala 292:{9,9}]
  wire [2:0] vCSR_2_frm = CSRFile_2_io_frm; // @[CSR.scala 270:{19,19}]
  wire [2:0] _GEN_14 = 2'h2 == io_frm_wid ? vCSR_2_frm : _GEN_13; // @[CSR.scala 292:{9,9}]
  wire [2:0] vCSR_3_frm = CSRFile_3_io_frm; // @[CSR.scala 270:{19,19}]
  CSRFile CSRFile ( // @[CSR.scala 270:45]
    .clock(CSRFile_clock),
    .reset(CSRFile_reset),
    .io_ctrl_inst(CSRFile_io_ctrl_inst),
    .io_ctrl_csr(CSRFile_io_ctrl_csr),
    .io_ctrl_isvec(CSRFile_io_ctrl_isvec),
    .io_in1(CSRFile_io_in1),
    .io_write(CSRFile_io_write),
    .io_wb_wxd_rd(CSRFile_io_wb_wxd_rd),
    .io_frm(CSRFile_io_frm),
    .io_CTA2csr_valid(CSRFile_io_CTA2csr_valid),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count(CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch(CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch(CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch(CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch
      )
  );
  CSRFile CSRFile_1 ( // @[CSR.scala 270:45]
    .clock(CSRFile_1_clock),
    .reset(CSRFile_1_reset),
    .io_ctrl_inst(CSRFile_1_io_ctrl_inst),
    .io_ctrl_csr(CSRFile_1_io_ctrl_csr),
    .io_ctrl_isvec(CSRFile_1_io_ctrl_isvec),
    .io_in1(CSRFile_1_io_in1),
    .io_write(CSRFile_1_io_write),
    .io_wb_wxd_rd(CSRFile_1_io_wb_wxd_rd),
    .io_frm(CSRFile_1_io_frm),
    .io_CTA2csr_valid(CSRFile_1_io_CTA2csr_valid),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count(CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch(CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch
      ),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch(CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch(
      CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch)
  );
  CSRFile CSRFile_2 ( // @[CSR.scala 270:45]
    .clock(CSRFile_2_clock),
    .reset(CSRFile_2_reset),
    .io_ctrl_inst(CSRFile_2_io_ctrl_inst),
    .io_ctrl_csr(CSRFile_2_io_ctrl_csr),
    .io_ctrl_isvec(CSRFile_2_io_ctrl_isvec),
    .io_in1(CSRFile_2_io_in1),
    .io_write(CSRFile_2_io_write),
    .io_wb_wxd_rd(CSRFile_2_io_wb_wxd_rd),
    .io_frm(CSRFile_2_io_frm),
    .io_CTA2csr_valid(CSRFile_2_io_CTA2csr_valid),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count(CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch(CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch
      ),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch(CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch(
      CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch)
  );
  CSRFile CSRFile_3 ( // @[CSR.scala 270:45]
    .clock(CSRFile_3_clock),
    .reset(CSRFile_3_reset),
    .io_ctrl_inst(CSRFile_3_io_ctrl_inst),
    .io_ctrl_csr(CSRFile_3_io_ctrl_csr),
    .io_ctrl_isvec(CSRFile_3_io_ctrl_isvec),
    .io_in1(CSRFile_3_io_in1),
    .io_write(CSRFile_3_io_write),
    .io_wb_wxd_rd(CSRFile_3_io_wb_wxd_rd),
    .io_frm(CSRFile_3_io_frm),
    .io_CTA2csr_valid(CSRFile_3_io_CTA2csr_valid),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count(CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch(CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch
      ),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch(CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch(
      CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch)
  );
  Queue_1 result ( // @[CSR.scala 280:20]
    .clock(result_clock),
    .reset(result_reset),
    .io_enq_ready(result_io_enq_ready),
    .io_enq_valid(result_io_enq_valid),
    .io_enq_bits_wb_wxd_rd(result_io_enq_bits_wb_wxd_rd),
    .io_enq_bits_wxd(result_io_enq_bits_wxd),
    .io_enq_bits_reg_idxw(result_io_enq_bits_reg_idxw),
    .io_enq_bits_warp_id(result_io_enq_bits_warp_id),
    .io_deq_ready(result_io_deq_ready),
    .io_deq_valid(result_io_deq_valid),
    .io_deq_bits_wb_wxd_rd(result_io_deq_bits_wb_wxd_rd),
    .io_deq_bits_wxd(result_io_deq_bits_wxd),
    .io_deq_bits_reg_idxw(result_io_deq_bits_reg_idxw),
    .io_deq_bits_warp_id(result_io_deq_bits_warp_id)
  );
  assign io_in_ready = result_io_enq_ready & ~io_CTA2csr_valid; // @[CSR.scala 283:36]
  assign io_out_valid = result_io_deq_valid; // @[CSR.scala 281:16]
  assign io_out_bits_wb_wxd_rd = result_io_deq_bits_wb_wxd_rd; // @[CSR.scala 281:16]
  assign io_out_bits_wxd = result_io_deq_bits_wxd; // @[CSR.scala 281:16]
  assign io_out_bits_reg_idxw = result_io_deq_bits_reg_idxw; // @[CSR.scala 281:16]
  assign io_out_bits_warp_id = result_io_deq_bits_warp_id; // @[CSR.scala 281:16]
  assign io_frm = 2'h3 == io_frm_wid ? vCSR_3_frm : _GEN_14; // @[CSR.scala 292:{9,9}]
  assign CSRFile_clock = clock;
  assign CSRFile_reset = reset;
  assign CSRFile_io_ctrl_inst = io_in_bits_ctrl_inst; // @[CSR.scala 270:19 272:11]
  assign CSRFile_io_ctrl_csr = io_in_bits_ctrl_csr; // @[CSR.scala 270:19 272:11]
  assign CSRFile_io_ctrl_isvec = io_in_bits_ctrl_isvec; // @[CSR.scala 270:19 272:11]
  assign CSRFile_io_in1 = io_in_bits_in1; // @[CSR.scala 270:19 274:10]
  assign CSRFile_io_write = 2'h0 == io_in_bits_ctrl_wid & _vCSR_write_T; // @[CSR.scala 273:12 278:{34,34}]
  assign CSRFile_io_CTA2csr_valid = 2'h0 == io_CTA2csr_bits_wid & io_CTA2csr_valid; // @[CSR.scala 275:20 279:{42,42}]
  assign CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count = io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:19 276:19]
  assign CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_1_clock = clock;
  assign CSRFile_1_reset = reset;
  assign CSRFile_1_io_ctrl_inst = io_in_bits_ctrl_inst; // @[CSR.scala 270:19 272:11]
  assign CSRFile_1_io_ctrl_csr = io_in_bits_ctrl_csr; // @[CSR.scala 270:19 272:11]
  assign CSRFile_1_io_ctrl_isvec = io_in_bits_ctrl_isvec; // @[CSR.scala 270:19 272:11]
  assign CSRFile_1_io_in1 = io_in_bits_in1; // @[CSR.scala 270:19 274:10]
  assign CSRFile_1_io_write = 2'h1 == io_in_bits_ctrl_wid & _vCSR_write_T; // @[CSR.scala 273:12 278:{34,34}]
  assign CSRFile_1_io_CTA2csr_valid = 2'h1 == io_CTA2csr_bits_wid & io_CTA2csr_valid; // @[CSR.scala 275:20 279:{42,42}]
  assign CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count = io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:19 276:19]
  assign CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_1_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_2_clock = clock;
  assign CSRFile_2_reset = reset;
  assign CSRFile_2_io_ctrl_inst = io_in_bits_ctrl_inst; // @[CSR.scala 270:19 272:11]
  assign CSRFile_2_io_ctrl_csr = io_in_bits_ctrl_csr; // @[CSR.scala 270:19 272:11]
  assign CSRFile_2_io_ctrl_isvec = io_in_bits_ctrl_isvec; // @[CSR.scala 270:19 272:11]
  assign CSRFile_2_io_in1 = io_in_bits_in1; // @[CSR.scala 270:19 274:10]
  assign CSRFile_2_io_write = 2'h2 == io_in_bits_ctrl_wid & _vCSR_write_T; // @[CSR.scala 273:12 278:{34,34}]
  assign CSRFile_2_io_CTA2csr_valid = 2'h2 == io_CTA2csr_bits_wid & io_CTA2csr_valid; // @[CSR.scala 275:20 279:{42,42}]
  assign CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count = io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:19 276:19]
  assign CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_2_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_3_clock = clock;
  assign CSRFile_3_reset = reset;
  assign CSRFile_3_io_ctrl_inst = io_in_bits_ctrl_inst; // @[CSR.scala 270:19 272:11]
  assign CSRFile_3_io_ctrl_csr = io_in_bits_ctrl_csr; // @[CSR.scala 270:19 272:11]
  assign CSRFile_3_io_ctrl_isvec = io_in_bits_ctrl_isvec; // @[CSR.scala 270:19 272:11]
  assign CSRFile_3_io_in1 = io_in_bits_in1; // @[CSR.scala 270:19 274:10]
  assign CSRFile_3_io_write = 2'h3 == io_in_bits_ctrl_wid & _vCSR_write_T; // @[CSR.scala 273:12 278:{34,34}]
  assign CSRFile_3_io_CTA2csr_valid = 2'h3 == io_CTA2csr_bits_wid & io_CTA2csr_valid; // @[CSR.scala 275:20 279:{42,42}]
  assign CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count = io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[CSR.scala 270:19 276:19]
  assign CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[CSR.scala 270:19 276:19]
  assign CSRFile_3_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[CSR.scala 270:19 276:19]
  assign result_clock = clock;
  assign result_reset = reset;
  assign result_io_enq_valid = io_in_valid; // @[CSR.scala 284:22]
  assign result_io_enq_bits_wb_wxd_rd = 2'h3 == io_in_bits_ctrl_wid ? vCSR_3_wb_wxd_rd : _GEN_10; // @[CSR.scala 288:{31,31}]
  assign result_io_enq_bits_wxd = io_in_bits_ctrl_wxd; // @[CSR.scala 287:25]
  assign result_io_enq_bits_reg_idxw = io_in_bits_ctrl_reg_idxw; // @[CSR.scala 286:30]
  assign result_io_enq_bits_warp_id = io_in_bits_ctrl_wid; // @[CSR.scala 289:29]
  assign result_io_deq_ready = io_out_ready; // @[CSR.scala 281:16]
endmodule
module pipe(
  input         clock,
  input         reset,
  output        io_icache_req_valid,
  output [31:0] io_icache_req_bits_addr,
  output [1:0]  io_icache_req_bits_warpid,
  input         io_icache_rsp_valid,
  input  [31:0] io_icache_rsp_bits_addr,
  input  [31:0] io_icache_rsp_bits_data,
  input  [1:0]  io_icache_rsp_bits_warpid,
  input  [1:0]  io_icache_rsp_bits_status,
  output        io_externalFlushPipe_valid,
  output [1:0]  io_externalFlushPipe_bits,
  input         io_dcache_req_ready,
  output        io_dcache_req_valid,
  output [1:0]  io_dcache_req_bits_instrId,
  output        io_dcache_req_bits_isWrite,
  output [21:0] io_dcache_req_bits_tag,
  output [4:0]  io_dcache_req_bits_setIdx,
  output        io_dcache_req_bits_perLaneAddr_0_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_0_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_1_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_1_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_2_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_2_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_3_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_3_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_4_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_4_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_5_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_5_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_6_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_6_blockOffset,
  output        io_dcache_req_bits_perLaneAddr_7_activeMask,
  output [2:0]  io_dcache_req_bits_perLaneAddr_7_blockOffset,
  output [31:0] io_dcache_req_bits_data_0,
  output [31:0] io_dcache_req_bits_data_1,
  output [31:0] io_dcache_req_bits_data_2,
  output [31:0] io_dcache_req_bits_data_3,
  output [31:0] io_dcache_req_bits_data_4,
  output [31:0] io_dcache_req_bits_data_5,
  output [31:0] io_dcache_req_bits_data_6,
  output [31:0] io_dcache_req_bits_data_7,
  output        io_dcache_rsp_ready,
  input         io_dcache_rsp_valid,
  input  [1:0]  io_dcache_rsp_bits_instrId,
  input  [31:0] io_dcache_rsp_bits_data_0,
  input  [31:0] io_dcache_rsp_bits_data_1,
  input  [31:0] io_dcache_rsp_bits_data_2,
  input  [31:0] io_dcache_rsp_bits_data_3,
  input  [31:0] io_dcache_rsp_bits_data_4,
  input  [31:0] io_dcache_rsp_bits_data_5,
  input  [31:0] io_dcache_rsp_bits_data_6,
  input  [31:0] io_dcache_rsp_bits_data_7,
  input         io_dcache_rsp_bits_activeMask_0,
  input         io_dcache_rsp_bits_activeMask_1,
  input         io_dcache_rsp_bits_activeMask_2,
  input         io_dcache_rsp_bits_activeMask_3,
  input         io_dcache_rsp_bits_activeMask_4,
  input         io_dcache_rsp_bits_activeMask_5,
  input         io_dcache_rsp_bits_activeMask_6,
  input         io_dcache_rsp_bits_activeMask_7,
  input         io_shared_req_ready,
  output        io_shared_req_valid,
  output [1:0]  io_shared_req_bits_instrId,
  output        io_shared_req_bits_isWrite,
  output [4:0]  io_shared_req_bits_setIdx,
  output        io_shared_req_bits_perLaneAddr_0_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_0_blockOffset,
  output        io_shared_req_bits_perLaneAddr_1_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_1_blockOffset,
  output        io_shared_req_bits_perLaneAddr_2_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_2_blockOffset,
  output        io_shared_req_bits_perLaneAddr_3_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_3_blockOffset,
  output        io_shared_req_bits_perLaneAddr_4_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_4_blockOffset,
  output        io_shared_req_bits_perLaneAddr_5_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_5_blockOffset,
  output        io_shared_req_bits_perLaneAddr_6_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_6_blockOffset,
  output        io_shared_req_bits_perLaneAddr_7_activeMask,
  output [2:0]  io_shared_req_bits_perLaneAddr_7_blockOffset,
  output [31:0] io_shared_req_bits_data_0,
  output [31:0] io_shared_req_bits_data_1,
  output [31:0] io_shared_req_bits_data_2,
  output [31:0] io_shared_req_bits_data_3,
  output [31:0] io_shared_req_bits_data_4,
  output [31:0] io_shared_req_bits_data_5,
  output [31:0] io_shared_req_bits_data_6,
  output [31:0] io_shared_req_bits_data_7,
  output        io_shared_rsp_ready,
  input         io_shared_rsp_valid,
  input  [1:0]  io_shared_rsp_bits_instrId,
  input  [31:0] io_shared_rsp_bits_data_0,
  input  [31:0] io_shared_rsp_bits_data_1,
  input  [31:0] io_shared_rsp_bits_data_2,
  input  [31:0] io_shared_rsp_bits_data_3,
  input  [31:0] io_shared_rsp_bits_data_4,
  input  [31:0] io_shared_rsp_bits_data_5,
  input  [31:0] io_shared_rsp_bits_data_6,
  input  [31:0] io_shared_rsp_bits_data_7,
  input         io_shared_rsp_bits_activeMask_0,
  input         io_shared_rsp_bits_activeMask_1,
  input         io_shared_rsp_bits_activeMask_2,
  input         io_shared_rsp_bits_activeMask_3,
  input         io_shared_rsp_bits_activeMask_4,
  input         io_shared_rsp_bits_activeMask_5,
  input         io_shared_rsp_bits_activeMask_6,
  input         io_shared_rsp_bits_activeMask_7,
  input         io_pc_reset,
  input         io_warpReq_valid,
  input  [2:0]  io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count,
  input  [9:0]  io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch,
  input  [12:0] io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch,
  input  [12:0] io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch,
  input  [4:0]  io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch,
  input  [12:0] io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch,
  input  [31:0] io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch,
  input  [1:0]  io_warpReq_bits_wid,
  output        io_warpRsp_valid,
  output [1:0]  io_warpRsp_bits_wid,
  output [1:0]  io_wg_id_lookup,
  input  [4:0]  io_wg_id_tag
);
  wire  warp_sche_clock; // @[pipe.scala 39:23]
  wire  warp_sche_reset; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_reset; // @[pipe.scala 39:23]
  wire  warp_sche_io_warpReq_ready; // @[pipe.scala 39:23]
  wire  warp_sche_io_warpReq_valid; // @[pipe.scala 39:23]
  wire [2:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count; // @[pipe.scala 39:23]
  wire [9:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[pipe.scala 39:23]
  wire [12:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[pipe.scala 39:23]
  wire [12:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[pipe.scala 39:23]
  wire [4:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[pipe.scala 39:23]
  wire [12:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[pipe.scala 39:23]
  wire [31:0] warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_warpReq_bits_wid; // @[pipe.scala 39:23]
  wire  warp_sche_io_warpRsp_valid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_warpRsp_bits_wid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_wg_id_lookup; // @[pipe.scala 39:23]
  wire [4:0] warp_sche_io_wg_id_tag; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_req_valid; // @[pipe.scala 39:23]
  wire [31:0] warp_sche_io_pc_req_bits_addr; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_pc_req_bits_warpid; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_rsp_valid; // @[pipe.scala 39:23]
  wire [31:0] warp_sche_io_pc_rsp_bits_addr; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_pc_rsp_bits_warpid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_pc_rsp_bits_status; // @[pipe.scala 39:23]
  wire  warp_sche_io_branch_ready; // @[pipe.scala 39:23]
  wire  warp_sche_io_branch_valid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_branch_bits_wid; // @[pipe.scala 39:23]
  wire  warp_sche_io_branch_bits_jump; // @[pipe.scala 39:23]
  wire [31:0] warp_sche_io_branch_bits_new_pc; // @[pipe.scala 39:23]
  wire  warp_sche_io_warp_control_ready; // @[pipe.scala 39:23]
  wire  warp_sche_io_warp_control_valid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_warp_control_bits_ctrl_wid; // @[pipe.scala 39:23]
  wire  warp_sche_io_warp_control_bits_ctrl_simt_stack_op; // @[pipe.scala 39:23]
  wire  warp_sche_io_warp_control_bits_ctrl_barrier; // @[pipe.scala 39:23]
  wire [3:0] warp_sche_io_scoreboard_busy; // @[pipe.scala 39:23]
  wire [3:0] warp_sche_io_exe_busy; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_ibuffer_ready_0; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_ibuffer_ready_1; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_ibuffer_ready_2; // @[pipe.scala 39:23]
  wire  warp_sche_io_pc_ibuffer_ready_3; // @[pipe.scala 39:23]
  wire [3:0] warp_sche_io_warp_ready; // @[pipe.scala 39:23]
  wire  warp_sche_io_flush_valid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_flush_bits; // @[pipe.scala 39:23]
  wire  warp_sche_io_flushCache_valid; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_flushCache_bits; // @[pipe.scala 39:23]
  wire  warp_sche_io_CTA2csr_valid; // @[pipe.scala 39:23]
  wire [2:0] warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[pipe.scala 39:23]
  wire [9:0] warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[pipe.scala 39:23]
  wire [12:0] warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[pipe.scala 39:23]
  wire [12:0] warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[pipe.scala 39:23]
  wire [4:0] warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[pipe.scala 39:23]
  wire [12:0] warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[pipe.scala 39:23]
  wire [1:0] warp_sche_io_CTA2csr_bits_wid; // @[pipe.scala 39:23]
  wire [31:0] control_io_inst; // @[pipe.scala 41:21]
  wire [31:0] control_io_pc; // @[pipe.scala 41:21]
  wire [1:0] control_io_wid; // @[pipe.scala 41:21]
  wire [31:0] control_io_control_inst; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_wid; // @[pipe.scala 41:21]
  wire  control_io_control_fp; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_branch; // @[pipe.scala 41:21]
  wire  control_io_control_simt_stack; // @[pipe.scala 41:21]
  wire  control_io_control_simt_stack_op; // @[pipe.scala 41:21]
  wire  control_io_control_barrier; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_csr; // @[pipe.scala 41:21]
  wire  control_io_control_reverse; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_sel_alu2; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_sel_alu1; // @[pipe.scala 41:21]
  wire  control_io_control_isvec; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_sel_alu3; // @[pipe.scala 41:21]
  wire  control_io_control_mask; // @[pipe.scala 41:21]
  wire [2:0] control_io_control_sel_imm; // @[pipe.scala 41:21]
  wire  control_io_control_mem_unsigned; // @[pipe.scala 41:21]
  wire [5:0] control_io_control_alu_fn; // @[pipe.scala 41:21]
  wire  control_io_control_mem; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_mem_cmd; // @[pipe.scala 41:21]
  wire [1:0] control_io_control_mop; // @[pipe.scala 41:21]
  wire [4:0] control_io_control_reg_idx1; // @[pipe.scala 41:21]
  wire [4:0] control_io_control_reg_idx2; // @[pipe.scala 41:21]
  wire [4:0] control_io_control_reg_idx3; // @[pipe.scala 41:21]
  wire [4:0] control_io_control_reg_idxw; // @[pipe.scala 41:21]
  wire  control_io_control_wfd; // @[pipe.scala 41:21]
  wire  control_io_control_fence; // @[pipe.scala 41:21]
  wire  control_io_control_sfu; // @[pipe.scala 41:21]
  wire  control_io_control_readmask; // @[pipe.scala 41:21]
  wire  control_io_control_writemask; // @[pipe.scala 41:21]
  wire  control_io_control_wxd; // @[pipe.scala 41:21]
  wire [31:0] control_io_control_pc; // @[pipe.scala 41:21]
  wire  operand_collector_clock; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_control_inst; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_control_wid; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_control_branch; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_control_sel_alu2; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_control_sel_alu1; // @[pipe.scala 42:31]
  wire  operand_collector_io_control_isvec; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_control_sel_alu3; // @[pipe.scala 42:31]
  wire  operand_collector_io_control_mask; // @[pipe.scala 42:31]
  wire [2:0] operand_collector_io_control_sel_imm; // @[pipe.scala 42:31]
  wire [4:0] operand_collector_io_control_reg_idx1; // @[pipe.scala 42:31]
  wire [4:0] operand_collector_io_control_reg_idx2; // @[pipe.scala 42:31]
  wire [4:0] operand_collector_io_control_reg_idx3; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_control_pc; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_0; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_1; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_2; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_3; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_4; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_5; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_6; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src1_7; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_0; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_1; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_2; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_3; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_4; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_5; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_6; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src2_7; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_0; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_1; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_2; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_3; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_4; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_5; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_6; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_alu_src3_7; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_0; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_1; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_2; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_3; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_4; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_5; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_6; // @[pipe.scala 42:31]
  wire  operand_collector_io_mask_7; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeScalarCtrl_valid; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeScalarCtrl_bits_wb_wxd_rd; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeScalarCtrl_bits_wxd; // @[pipe.scala 42:31]
  wire [4:0] operand_collector_io_writeScalarCtrl_bits_reg_idxw; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_writeScalarCtrl_bits_warp_id; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_valid; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_0; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_1; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_2; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_3; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_4; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_5; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_6; // @[pipe.scala 42:31]
  wire [31:0] operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_7; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_0; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_1; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_2; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_3; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_4; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_5; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_6; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd_mask_7; // @[pipe.scala 42:31]
  wire  operand_collector_io_writeVecCtrl_bits_wfd; // @[pipe.scala 42:31]
  wire [4:0] operand_collector_io_writeVecCtrl_bits_reg_idxw; // @[pipe.scala 42:31]
  wire [1:0] operand_collector_io_writeVecCtrl_bits_warp_id; // @[pipe.scala 42:31]
  wire  issue_io_in_ready; // @[pipe.scala 43:19]
  wire  issue_io_in_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in1_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in2_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_in3_7; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_0; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_1; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_2; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_3; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_4; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_5; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_6; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_mask_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_ctrl_inst; // @[pipe.scala 43:19]
  wire [1:0] issue_io_in_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_fp; // @[pipe.scala 43:19]
  wire [1:0] issue_io_in_bits_ctrl_branch; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_simt_stack; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_simt_stack_op; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_barrier; // @[pipe.scala 43:19]
  wire [1:0] issue_io_in_bits_ctrl_csr; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_reverse; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_isvec; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_mem_unsigned; // @[pipe.scala 43:19]
  wire [5:0] issue_io_in_bits_ctrl_alu_fn; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_mem; // @[pipe.scala 43:19]
  wire [1:0] issue_io_in_bits_ctrl_mem_cmd; // @[pipe.scala 43:19]
  wire [1:0] issue_io_in_bits_ctrl_mop; // @[pipe.scala 43:19]
  wire [4:0] issue_io_in_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_wfd; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_fence; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_sfu; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_readmask; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_writemask; // @[pipe.scala 43:19]
  wire  issue_io_in_bits_ctrl_wxd; // @[pipe.scala 43:19]
  wire [31:0] issue_io_in_bits_ctrl_pc; // @[pipe.scala 43:19]
  wire  issue_io_out_sALU_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_sALU_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_sALU_bits_in1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_sALU_bits_in2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_sALU_bits_in3; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_sALU_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_sALU_bits_ctrl_branch; // @[pipe.scala 43:19]
  wire [5:0] issue_io_out_sALU_bits_ctrl_alu_fn; // @[pipe.scala 43:19]
  wire [4:0] issue_io_out_sALU_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_out_sALU_bits_ctrl_wxd; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in1_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in2_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vALU_bits_in3_7; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_0; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_1; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_2; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_3; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_4; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_5; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_6; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_mask_7; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_vALU_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_ctrl_simt_stack; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_ctrl_reverse; // @[pipe.scala 43:19]
  wire [5:0] issue_io_out_vALU_bits_ctrl_alu_fn; // @[pipe.scala 43:19]
  wire [4:0] issue_io_out_vALU_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_ctrl_wfd; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_ctrl_readmask; // @[pipe.scala 43:19]
  wire  issue_io_out_vALU_bits_ctrl_writemask; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in1_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in2_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_vFPU_bits_in3_7; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_0; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_1; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_2; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_3; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_4; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_5; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_6; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_mask_7; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_vFPU_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_ctrl_reverse; // @[pipe.scala 43:19]
  wire [5:0] issue_io_out_vFPU_bits_ctrl_alu_fn; // @[pipe.scala 43:19]
  wire [4:0] issue_io_out_vFPU_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_ctrl_wfd; // @[pipe.scala 43:19]
  wire  issue_io_out_vFPU_bits_ctrl_wxd; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in1_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in2_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_in3_7; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_0; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_1; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_2; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_3; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_4; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_5; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_6; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_mask_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_ctrl_inst; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_LSU_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_fp; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_LSU_bits_ctrl_branch; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_simt_stack; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_simt_stack_op; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_barrier; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_LSU_bits_ctrl_csr; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_reverse; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_isvec; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_mem_unsigned; // @[pipe.scala 43:19]
  wire [5:0] issue_io_out_LSU_bits_ctrl_alu_fn; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_mem; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_LSU_bits_ctrl_mem_cmd; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_LSU_bits_ctrl_mop; // @[pipe.scala 43:19]
  wire [4:0] issue_io_out_LSU_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_wfd; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_fence; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_sfu; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_readmask; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_writemask; // @[pipe.scala 43:19]
  wire  issue_io_out_LSU_bits_ctrl_wxd; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_LSU_bits_ctrl_pc; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in1_7; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_0; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_1; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_2; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_3; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_4; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_5; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_6; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SFU_bits_in2_7; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_0; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_1; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_2; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_3; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_4; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_5; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_6; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_mask_7; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_SFU_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_ctrl_fp; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_ctrl_reverse; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_ctrl_isvec; // @[pipe.scala 43:19]
  wire [5:0] issue_io_out_SFU_bits_ctrl_alu_fn; // @[pipe.scala 43:19]
  wire [4:0] issue_io_out_SFU_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_ctrl_wfd; // @[pipe.scala 43:19]
  wire  issue_io_out_SFU_bits_ctrl_wxd; // @[pipe.scala 43:19]
  wire  issue_io_out_SIMT_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_SIMT_valid; // @[pipe.scala 43:19]
  wire  issue_io_out_SIMT_bits_opcode; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_SIMT_bits_wid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_SIMT_bits_PC_branch; // @[pipe.scala 43:19]
  wire [7:0] issue_io_out_SIMT_bits_mask_init; // @[pipe.scala 43:19]
  wire  issue_io_out_warpscheduler_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_warpscheduler_valid; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_warpscheduler_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire  issue_io_out_warpscheduler_bits_ctrl_simt_stack_op; // @[pipe.scala 43:19]
  wire  issue_io_out_warpscheduler_bits_ctrl_barrier; // @[pipe.scala 43:19]
  wire  issue_io_out_CSR_ready; // @[pipe.scala 43:19]
  wire  issue_io_out_CSR_valid; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_CSR_bits_ctrl_inst; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_CSR_bits_ctrl_wid; // @[pipe.scala 43:19]
  wire [1:0] issue_io_out_CSR_bits_ctrl_csr; // @[pipe.scala 43:19]
  wire  issue_io_out_CSR_bits_ctrl_isvec; // @[pipe.scala 43:19]
  wire [4:0] issue_io_out_CSR_bits_ctrl_reg_idxw; // @[pipe.scala 43:19]
  wire  issue_io_out_CSR_bits_ctrl_wxd; // @[pipe.scala 43:19]
  wire [31:0] issue_io_out_CSR_bits_in1; // @[pipe.scala 43:19]
  wire  alu_clock; // @[pipe.scala 44:17]
  wire  alu_reset; // @[pipe.scala 44:17]
  wire  alu_io_in_ready; // @[pipe.scala 44:17]
  wire  alu_io_in_valid; // @[pipe.scala 44:17]
  wire [31:0] alu_io_in_bits_in1; // @[pipe.scala 44:17]
  wire [31:0] alu_io_in_bits_in2; // @[pipe.scala 44:17]
  wire [31:0] alu_io_in_bits_in3; // @[pipe.scala 44:17]
  wire [1:0] alu_io_in_bits_ctrl_wid; // @[pipe.scala 44:17]
  wire [1:0] alu_io_in_bits_ctrl_branch; // @[pipe.scala 44:17]
  wire [5:0] alu_io_in_bits_ctrl_alu_fn; // @[pipe.scala 44:17]
  wire [4:0] alu_io_in_bits_ctrl_reg_idxw; // @[pipe.scala 44:17]
  wire  alu_io_in_bits_ctrl_wxd; // @[pipe.scala 44:17]
  wire  alu_io_out_valid; // @[pipe.scala 44:17]
  wire [31:0] alu_io_out_bits_wb_wxd_rd; // @[pipe.scala 44:17]
  wire  alu_io_out_bits_wxd; // @[pipe.scala 44:17]
  wire [4:0] alu_io_out_bits_reg_idxw; // @[pipe.scala 44:17]
  wire [1:0] alu_io_out_bits_warp_id; // @[pipe.scala 44:17]
  wire  alu_io_out2br_ready; // @[pipe.scala 44:17]
  wire  alu_io_out2br_valid; // @[pipe.scala 44:17]
  wire [1:0] alu_io_out2br_bits_wid; // @[pipe.scala 44:17]
  wire  alu_io_out2br_bits_jump; // @[pipe.scala 44:17]
  wire [31:0] alu_io_out2br_bits_new_pc; // @[pipe.scala 44:17]
  wire  valu_clock; // @[pipe.scala 45:18]
  wire  valu_reset; // @[pipe.scala 45:18]
  wire  valu_io_in_ready; // @[pipe.scala 45:18]
  wire  valu_io_in_valid; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_0; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_1; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_2; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_3; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_4; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_5; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_6; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in1_7; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_0; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_1; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_2; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_3; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_4; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_5; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_6; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in2_7; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_0; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_1; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_2; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_3; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_4; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_5; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_6; // @[pipe.scala 45:18]
  wire [31:0] valu_io_in_bits_in3_7; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_0; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_1; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_2; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_3; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_4; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_5; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_6; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_mask_7; // @[pipe.scala 45:18]
  wire [1:0] valu_io_in_bits_ctrl_wid; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_ctrl_simt_stack; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_ctrl_reverse; // @[pipe.scala 45:18]
  wire [5:0] valu_io_in_bits_ctrl_alu_fn; // @[pipe.scala 45:18]
  wire [4:0] valu_io_in_bits_ctrl_reg_idxw; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_ctrl_wfd; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_ctrl_readmask; // @[pipe.scala 45:18]
  wire  valu_io_in_bits_ctrl_writemask; // @[pipe.scala 45:18]
  wire  valu_io_out_valid; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_0; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_1; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_2; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_3; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_4; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_5; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_6; // @[pipe.scala 45:18]
  wire [31:0] valu_io_out_bits_wb_wfd_rd_7; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_0; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_1; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_2; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_3; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_4; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_5; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_6; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd_mask_7; // @[pipe.scala 45:18]
  wire  valu_io_out_bits_wfd; // @[pipe.scala 45:18]
  wire [4:0] valu_io_out_bits_reg_idxw; // @[pipe.scala 45:18]
  wire [1:0] valu_io_out_bits_warp_id; // @[pipe.scala 45:18]
  wire  valu_io_out2simt_stack_ready; // @[pipe.scala 45:18]
  wire  valu_io_out2simt_stack_valid; // @[pipe.scala 45:18]
  wire [7:0] valu_io_out2simt_stack_bits_if_mask; // @[pipe.scala 45:18]
  wire [1:0] valu_io_out2simt_stack_bits_wid; // @[pipe.scala 45:18]
  wire  fpu_clock; // @[pipe.scala 46:17]
  wire  fpu_reset; // @[pipe.scala 46:17]
  wire  fpu_io_in_ready; // @[pipe.scala 46:17]
  wire  fpu_io_in_valid; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_0; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_1; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_2; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_3; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_4; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_5; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_6; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in1_7; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_0; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_1; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_2; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_3; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_4; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_5; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_6; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in2_7; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_0; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_1; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_2; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_3; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_4; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_5; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_6; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_in_bits_in3_7; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_0; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_1; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_2; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_3; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_4; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_5; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_6; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_mask_7; // @[pipe.scala 46:17]
  wire [1:0] fpu_io_in_bits_ctrl_wid; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_ctrl_reverse; // @[pipe.scala 46:17]
  wire [5:0] fpu_io_in_bits_ctrl_alu_fn; // @[pipe.scala 46:17]
  wire [4:0] fpu_io_in_bits_ctrl_reg_idxw; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_ctrl_wfd; // @[pipe.scala 46:17]
  wire  fpu_io_in_bits_ctrl_wxd; // @[pipe.scala 46:17]
  wire [2:0] fpu_io_rm; // @[pipe.scala 46:17]
  wire  fpu_io_out_x_ready; // @[pipe.scala 46:17]
  wire  fpu_io_out_x_valid; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 46:17]
  wire  fpu_io_out_x_bits_wxd; // @[pipe.scala 46:17]
  wire [4:0] fpu_io_out_x_bits_reg_idxw; // @[pipe.scala 46:17]
  wire [1:0] fpu_io_out_x_bits_warp_id; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_ready; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_valid; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 46:17]
  wire [31:0] fpu_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_0; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_1; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_2; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_3; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_4; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_5; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_6; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd_mask_7; // @[pipe.scala 46:17]
  wire  fpu_io_out_v_bits_wfd; // @[pipe.scala 46:17]
  wire [4:0] fpu_io_out_v_bits_reg_idxw; // @[pipe.scala 46:17]
  wire [1:0] fpu_io_out_v_bits_warp_id; // @[pipe.scala 46:17]
  wire  lsu_clock; // @[pipe.scala 47:17]
  wire  lsu_reset; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_ready; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_valid; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in1_7; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in2_7; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_in3_7; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_0; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_1; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_2; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_3; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_4; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_5; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_6; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_mask_7; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_ctrl_inst; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_lsu_req_bits_ctrl_wid; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_fp; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_lsu_req_bits_ctrl_branch; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_simt_stack; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_simt_stack_op; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_barrier; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_lsu_req_bits_ctrl_csr; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_reverse; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_isvec; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_mem_unsigned; // @[pipe.scala 47:17]
  wire [5:0] lsu_io_lsu_req_bits_ctrl_alu_fn; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_mem; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_lsu_req_bits_ctrl_mem_cmd; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_lsu_req_bits_ctrl_mop; // @[pipe.scala 47:17]
  wire [4:0] lsu_io_lsu_req_bits_ctrl_reg_idxw; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_wfd; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_fence; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_sfu; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_readmask; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_writemask; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_req_bits_ctrl_wxd; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_req_bits_ctrl_pc; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_ready; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_valid; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_dcache_rsp_bits_instrId; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_rsp_bits_data_7; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_0; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_1; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_2; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_3; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_4; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_5; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_6; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_rsp_bits_activeMask_7; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_ready; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_valid; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_lsu_rsp_bits_tag_warp_id; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_wfd; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_wxd; // @[pipe.scala 47:17]
  wire [4:0] lsu_io_lsu_rsp_bits_tag_reg_idxw; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_0; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_1; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_2; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_3; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_4; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_5; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_6; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_mask_7; // @[pipe.scala 47:17]
  wire  lsu_io_lsu_rsp_bits_tag_isWrite; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_lsu_rsp_bits_data_7; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_ready; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_valid; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_dcache_req_bits_instrId; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_isWrite; // @[pipe.scala 47:17]
  wire [21:0] lsu_io_dcache_req_bits_tag; // @[pipe.scala 47:17]
  wire [4:0] lsu_io_dcache_req_bits_setIdx; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_0_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_0_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_1_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_1_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_2_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_2_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_3_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_3_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_4_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_4_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_5_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_5_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_6_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_6_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_dcache_req_bits_perLaneAddr_7_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_dcache_req_bits_perLaneAddr_7_blockOffset; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_dcache_req_bits_data_7; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_ready; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_valid; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_shared_req_bits_instrId; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_isWrite; // @[pipe.scala 47:17]
  wire [4:0] lsu_io_shared_req_bits_setIdx; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_0_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_0_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_1_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_1_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_2_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_2_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_3_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_3_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_4_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_4_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_5_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_5_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_6_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_6_blockOffset; // @[pipe.scala 47:17]
  wire  lsu_io_shared_req_bits_perLaneAddr_7_activeMask; // @[pipe.scala 47:17]
  wire [2:0] lsu_io_shared_req_bits_perLaneAddr_7_blockOffset; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_req_bits_data_7; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_ready; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_valid; // @[pipe.scala 47:17]
  wire [1:0] lsu_io_shared_rsp_bits_instrId; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_0; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_1; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_2; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_3; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_4; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_5; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_6; // @[pipe.scala 47:17]
  wire [31:0] lsu_io_shared_rsp_bits_data_7; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_0; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_1; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_2; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_3; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_4; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_5; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_6; // @[pipe.scala 47:17]
  wire  lsu_io_shared_rsp_bits_activeMask_7; // @[pipe.scala 47:17]
  wire [3:0] lsu_io_fence_end; // @[pipe.scala 47:17]
  wire  sfu_clock; // @[pipe.scala 48:17]
  wire  sfu_reset; // @[pipe.scala 48:17]
  wire  sfu_io_in_ready; // @[pipe.scala 48:17]
  wire  sfu_io_in_valid; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_0; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_1; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_2; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_3; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_4; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_5; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_6; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in1_7; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_0; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_1; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_2; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_3; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_4; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_5; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_6; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_in_bits_in2_7; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_0; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_1; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_2; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_3; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_4; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_5; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_6; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_mask_7; // @[pipe.scala 48:17]
  wire [1:0] sfu_io_in_bits_ctrl_wid; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_ctrl_fp; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_ctrl_reverse; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_ctrl_isvec; // @[pipe.scala 48:17]
  wire [5:0] sfu_io_in_bits_ctrl_alu_fn; // @[pipe.scala 48:17]
  wire [4:0] sfu_io_in_bits_ctrl_reg_idxw; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_ctrl_wfd; // @[pipe.scala 48:17]
  wire  sfu_io_in_bits_ctrl_wxd; // @[pipe.scala 48:17]
  wire [2:0] sfu_io_rm; // @[pipe.scala 48:17]
  wire  sfu_io_out_x_ready; // @[pipe.scala 48:17]
  wire  sfu_io_out_x_valid; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 48:17]
  wire  sfu_io_out_x_bits_wxd; // @[pipe.scala 48:17]
  wire [4:0] sfu_io_out_x_bits_reg_idxw; // @[pipe.scala 48:17]
  wire [1:0] sfu_io_out_x_bits_warp_id; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_ready; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_valid; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 48:17]
  wire [31:0] sfu_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_0; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_1; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_2; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_3; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_4; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_5; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_6; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd_mask_7; // @[pipe.scala 48:17]
  wire  sfu_io_out_v_bits_wfd; // @[pipe.scala 48:17]
  wire [4:0] sfu_io_out_v_bits_reg_idxw; // @[pipe.scala 48:17]
  wire [1:0] sfu_io_out_v_bits_warp_id; // @[pipe.scala 48:17]
  wire  lsu2wb_io_lsu_rsp_ready; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_valid; // @[pipe.scala 49:20]
  wire [1:0] lsu2wb_io_lsu_rsp_bits_tag_warp_id; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_wfd; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_wxd; // @[pipe.scala 49:20]
  wire [4:0] lsu2wb_io_lsu_rsp_bits_tag_reg_idxw; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_0; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_1; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_2; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_3; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_4; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_5; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_6; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_mask_7; // @[pipe.scala 49:20]
  wire  lsu2wb_io_lsu_rsp_bits_tag_isWrite; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_0; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_1; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_2; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_3; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_4; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_5; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_6; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_lsu_rsp_bits_data_7; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_x_ready; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_x_valid; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_x_bits_wxd; // @[pipe.scala 49:20]
  wire [4:0] lsu2wb_io_out_x_bits_reg_idxw; // @[pipe.scala 49:20]
  wire [1:0] lsu2wb_io_out_x_bits_warp_id; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_ready; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_valid; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 49:20]
  wire [31:0] lsu2wb_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_0; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_1; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_2; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_3; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_4; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_5; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_6; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd_mask_7; // @[pipe.scala 49:20]
  wire  lsu2wb_io_out_v_bits_wfd; // @[pipe.scala 49:20]
  wire [4:0] lsu2wb_io_out_v_bits_reg_idxw; // @[pipe.scala 49:20]
  wire [1:0] lsu2wb_io_out_v_bits_warp_id; // @[pipe.scala 49:20]
  wire  wb_io_out_v_ready; // @[pipe.scala 50:16]
  wire  wb_io_out_v_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_0; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_1; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_2; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_3; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_4; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_5; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_6; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd_mask_7; // @[pipe.scala 50:16]
  wire  wb_io_out_v_bits_wfd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_out_v_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_out_v_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_out_x_ready; // @[pipe.scala 50:16]
  wire  wb_io_out_x_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 50:16]
  wire  wb_io_out_x_bits_wxd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_out_x_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_out_x_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_x_0_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_x_0_bits_wb_wxd_rd; // @[pipe.scala 50:16]
  wire  wb_io_in_x_0_bits_wxd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_x_0_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_x_0_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_x_1_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_x_1_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_x_1_bits_wb_wxd_rd; // @[pipe.scala 50:16]
  wire  wb_io_in_x_1_bits_wxd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_x_1_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_x_1_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_x_2_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_x_2_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_x_2_bits_wb_wxd_rd; // @[pipe.scala 50:16]
  wire  wb_io_in_x_2_bits_wxd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_x_2_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_x_2_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_x_3_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_x_3_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_x_3_bits_wb_wxd_rd; // @[pipe.scala 50:16]
  wire  wb_io_in_x_3_bits_wxd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_x_3_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_x_3_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_x_4_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_x_4_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_x_4_bits_wb_wxd_rd; // @[pipe.scala 50:16]
  wire  wb_io_in_x_4_bits_wxd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_x_4_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_x_4_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_0; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_1; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_2; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_3; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_4; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_5; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_6; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_0_bits_wb_wfd_rd_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_0; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_1; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_2; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_3; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_4; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_5; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_6; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd_mask_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_0_bits_wfd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_v_0_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_v_0_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_0; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_1; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_2; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_3; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_4; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_5; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_6; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_1_bits_wb_wfd_rd_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_0; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_1; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_2; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_3; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_4; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_5; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_6; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd_mask_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_1_bits_wfd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_v_1_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_v_1_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_0; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_1; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_2; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_3; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_4; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_5; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_6; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_2_bits_wb_wfd_rd_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_0; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_1; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_2; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_3; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_4; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_5; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_6; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd_mask_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_2_bits_wfd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_v_2_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_v_2_bits_warp_id; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_ready; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_valid; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_0; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_1; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_2; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_3; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_4; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_5; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_6; // @[pipe.scala 50:16]
  wire [31:0] wb_io_in_v_3_bits_wb_wfd_rd_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_0; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_1; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_2; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_3; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_4; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_5; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_6; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd_mask_7; // @[pipe.scala 50:16]
  wire  wb_io_in_v_3_bits_wfd; // @[pipe.scala 50:16]
  wire [4:0] wb_io_in_v_3_bits_reg_idxw; // @[pipe.scala 50:16]
  wire [1:0] wb_io_in_v_3_bits_warp_id; // @[pipe.scala 50:16]
  wire  Scoreboard_clock; // @[pipe.scala 52:47]
  wire  Scoreboard_reset; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_io_ibuffer_if_ctrl_sel_alu2; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_io_ibuffer_if_ctrl_sel_alu1; // @[pipe.scala 52:47]
  wire  Scoreboard_io_ibuffer_if_ctrl_isvec; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_io_ibuffer_if_ctrl_sel_alu3; // @[pipe.scala 52:47]
  wire  Scoreboard_io_ibuffer_if_ctrl_mask; // @[pipe.scala 52:47]
  wire  Scoreboard_io_ibuffer_if_ctrl_mem; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_io_ibuffer_if_ctrl_reg_idx1; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_io_ibuffer_if_ctrl_reg_idx2; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_io_ibuffer_if_ctrl_reg_idx3; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_io_if_ctrl_branch; // @[pipe.scala 52:47]
  wire  Scoreboard_io_if_ctrl_barrier; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_io_if_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_io_if_ctrl_wfd; // @[pipe.scala 52:47]
  wire  Scoreboard_io_if_ctrl_fence; // @[pipe.scala 52:47]
  wire  Scoreboard_io_if_ctrl_wxd; // @[pipe.scala 52:47]
  wire  Scoreboard_io_wb_v_ctrl_wfd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_io_wb_v_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_io_wb_x_ctrl_wxd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_io_wb_x_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_io_if_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_io_br_ctrl; // @[pipe.scala 52:47]
  wire  Scoreboard_io_fence_end; // @[pipe.scala 52:47]
  wire  Scoreboard_io_wb_v_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_io_wb_x_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_io_delay; // @[pipe.scala 52:47]
  wire  Scoreboard_1_clock; // @[pipe.scala 52:47]
  wire  Scoreboard_1_reset; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_1_io_ibuffer_if_ctrl_sel_alu2; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_1_io_ibuffer_if_ctrl_sel_alu1; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_ibuffer_if_ctrl_isvec; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_1_io_ibuffer_if_ctrl_sel_alu3; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_ibuffer_if_ctrl_mask; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_ibuffer_if_ctrl_mem; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_1_io_ibuffer_if_ctrl_reg_idx1; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_1_io_ibuffer_if_ctrl_reg_idx2; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_1_io_ibuffer_if_ctrl_reg_idx3; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_1_io_if_ctrl_branch; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_if_ctrl_barrier; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_1_io_if_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_if_ctrl_wfd; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_if_ctrl_fence; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_if_ctrl_wxd; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_wb_v_ctrl_wfd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_1_io_wb_v_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_wb_x_ctrl_wxd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_1_io_wb_x_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_if_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_br_ctrl; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_fence_end; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_wb_v_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_wb_x_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_1_io_delay; // @[pipe.scala 52:47]
  wire  Scoreboard_2_clock; // @[pipe.scala 52:47]
  wire  Scoreboard_2_reset; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_2_io_ibuffer_if_ctrl_sel_alu2; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_2_io_ibuffer_if_ctrl_sel_alu1; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_ibuffer_if_ctrl_isvec; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_2_io_ibuffer_if_ctrl_sel_alu3; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_ibuffer_if_ctrl_mask; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_ibuffer_if_ctrl_mem; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_2_io_ibuffer_if_ctrl_reg_idx1; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_2_io_ibuffer_if_ctrl_reg_idx2; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_2_io_ibuffer_if_ctrl_reg_idx3; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_2_io_if_ctrl_branch; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_if_ctrl_barrier; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_2_io_if_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_if_ctrl_wfd; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_if_ctrl_fence; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_if_ctrl_wxd; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_wb_v_ctrl_wfd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_2_io_wb_v_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_wb_x_ctrl_wxd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_2_io_wb_x_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_if_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_br_ctrl; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_fence_end; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_wb_v_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_wb_x_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_2_io_delay; // @[pipe.scala 52:47]
  wire  Scoreboard_3_clock; // @[pipe.scala 52:47]
  wire  Scoreboard_3_reset; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_3_io_ibuffer_if_ctrl_sel_alu2; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_3_io_ibuffer_if_ctrl_sel_alu1; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_ibuffer_if_ctrl_isvec; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_3_io_ibuffer_if_ctrl_sel_alu3; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_ibuffer_if_ctrl_mask; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_ibuffer_if_ctrl_mem; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_3_io_ibuffer_if_ctrl_reg_idx1; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_3_io_ibuffer_if_ctrl_reg_idx2; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_3_io_ibuffer_if_ctrl_reg_idx3; // @[pipe.scala 52:47]
  wire [1:0] Scoreboard_3_io_if_ctrl_branch; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_if_ctrl_barrier; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_3_io_if_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_if_ctrl_wfd; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_if_ctrl_fence; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_if_ctrl_wxd; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_wb_v_ctrl_wfd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_3_io_wb_v_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_wb_x_ctrl_wxd; // @[pipe.scala 52:47]
  wire [4:0] Scoreboard_3_io_wb_x_ctrl_reg_idxw; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_if_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_br_ctrl; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_fence_end; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_wb_v_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_wb_x_fire; // @[pipe.scala 52:47]
  wire  Scoreboard_3_io_delay; // @[pipe.scala 52:47]
  wire  ibuffer_clock; // @[pipe.scala 53:21]
  wire  ibuffer_reset; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_ready; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_valid; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_in_bits_inst; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_wid; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_fp; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_branch; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_simt_stack; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_simt_stack_op; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_barrier; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_csr; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_reverse; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_sel_alu2; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_sel_alu1; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_isvec; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_sel_alu3; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_mask; // @[pipe.scala 53:21]
  wire [2:0] ibuffer_io_in_bits_sel_imm; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_mem_unsigned; // @[pipe.scala 53:21]
  wire [5:0] ibuffer_io_in_bits_alu_fn; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_mem; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_mem_cmd; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_in_bits_mop; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_in_bits_reg_idx1; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_in_bits_reg_idx2; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_in_bits_reg_idx3; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_in_bits_reg_idxw; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_wfd; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_fence; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_sfu; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_readmask; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_writemask; // @[pipe.scala 53:21]
  wire  ibuffer_io_in_bits_wxd; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_in_bits_pc; // @[pipe.scala 53:21]
  wire  ibuffer_io_flush_valid; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_flush_bits; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_ready; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_valid; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_0_bits_inst; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_wid; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_fp; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_branch; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_simt_stack; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_simt_stack_op; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_barrier; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_csr; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_reverse; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_sel_alu2; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_sel_alu1; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_isvec; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_sel_alu3; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_mask; // @[pipe.scala 53:21]
  wire [2:0] ibuffer_io_out_0_bits_sel_imm; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_mem_unsigned; // @[pipe.scala 53:21]
  wire [5:0] ibuffer_io_out_0_bits_alu_fn; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_mem; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_mem_cmd; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_0_bits_mop; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_0_bits_reg_idx1; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_0_bits_reg_idx2; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_0_bits_reg_idx3; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_0_bits_reg_idxw; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_wfd; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_fence; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_sfu; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_readmask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_writemask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_0_bits_wxd; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_0_bits_pc; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_ready; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_valid; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_1_bits_inst; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_wid; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_fp; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_branch; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_simt_stack; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_simt_stack_op; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_barrier; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_csr; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_reverse; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_sel_alu2; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_sel_alu1; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_isvec; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_sel_alu3; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_mask; // @[pipe.scala 53:21]
  wire [2:0] ibuffer_io_out_1_bits_sel_imm; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_mem_unsigned; // @[pipe.scala 53:21]
  wire [5:0] ibuffer_io_out_1_bits_alu_fn; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_mem; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_mem_cmd; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_1_bits_mop; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_1_bits_reg_idx1; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_1_bits_reg_idx2; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_1_bits_reg_idx3; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_1_bits_reg_idxw; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_wfd; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_fence; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_sfu; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_readmask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_writemask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_1_bits_wxd; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_1_bits_pc; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_ready; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_valid; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_2_bits_inst; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_wid; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_fp; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_branch; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_simt_stack; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_simt_stack_op; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_barrier; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_csr; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_reverse; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_sel_alu2; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_sel_alu1; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_isvec; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_sel_alu3; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_mask; // @[pipe.scala 53:21]
  wire [2:0] ibuffer_io_out_2_bits_sel_imm; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_mem_unsigned; // @[pipe.scala 53:21]
  wire [5:0] ibuffer_io_out_2_bits_alu_fn; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_mem; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_mem_cmd; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_2_bits_mop; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_2_bits_reg_idx1; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_2_bits_reg_idx2; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_2_bits_reg_idx3; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_2_bits_reg_idxw; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_wfd; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_fence; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_sfu; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_readmask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_writemask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_2_bits_wxd; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_2_bits_pc; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_ready; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_valid; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_3_bits_inst; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_wid; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_fp; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_branch; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_simt_stack; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_simt_stack_op; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_barrier; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_csr; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_reverse; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_sel_alu2; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_sel_alu1; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_isvec; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_sel_alu3; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_mask; // @[pipe.scala 53:21]
  wire [2:0] ibuffer_io_out_3_bits_sel_imm; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_mem_unsigned; // @[pipe.scala 53:21]
  wire [5:0] ibuffer_io_out_3_bits_alu_fn; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_mem; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_mem_cmd; // @[pipe.scala 53:21]
  wire [1:0] ibuffer_io_out_3_bits_mop; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_3_bits_reg_idx1; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_3_bits_reg_idx2; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_3_bits_reg_idx3; // @[pipe.scala 53:21]
  wire [4:0] ibuffer_io_out_3_bits_reg_idxw; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_wfd; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_fence; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_sfu; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_readmask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_writemask; // @[pipe.scala 53:21]
  wire  ibuffer_io_out_3_bits_wxd; // @[pipe.scala 53:21]
  wire [31:0] ibuffer_io_out_3_bits_pc; // @[pipe.scala 53:21]
  wire  ibuffer_io_ibuffer_ready_0; // @[pipe.scala 53:21]
  wire  ibuffer_io_ibuffer_ready_1; // @[pipe.scala 53:21]
  wire  ibuffer_io_ibuffer_ready_2; // @[pipe.scala 53:21]
  wire  ibuffer_io_ibuffer_ready_3; // @[pipe.scala 53:21]
  wire  ibuffer2issue_clock; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_ready; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_valid; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_0_bits_inst; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_wid; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_fp; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_branch; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_simt_stack; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_simt_stack_op; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_barrier; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_csr; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_reverse; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_sel_alu2; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_sel_alu1; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_isvec; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_sel_alu3; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_mask; // @[pipe.scala 54:27]
  wire [2:0] ibuffer2issue_io_in_0_bits_sel_imm; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_mem_unsigned; // @[pipe.scala 54:27]
  wire [5:0] ibuffer2issue_io_in_0_bits_alu_fn; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_mem; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_mem_cmd; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_0_bits_mop; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_0_bits_reg_idx1; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_0_bits_reg_idx2; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_0_bits_reg_idx3; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_0_bits_reg_idxw; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_wfd; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_fence; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_sfu; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_readmask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_writemask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_0_bits_wxd; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_0_bits_pc; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_ready; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_valid; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_1_bits_inst; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_wid; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_fp; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_branch; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_simt_stack; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_simt_stack_op; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_barrier; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_csr; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_reverse; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_sel_alu2; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_sel_alu1; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_isvec; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_sel_alu3; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_mask; // @[pipe.scala 54:27]
  wire [2:0] ibuffer2issue_io_in_1_bits_sel_imm; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_mem_unsigned; // @[pipe.scala 54:27]
  wire [5:0] ibuffer2issue_io_in_1_bits_alu_fn; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_mem; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_mem_cmd; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_1_bits_mop; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_1_bits_reg_idx1; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_1_bits_reg_idx2; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_1_bits_reg_idx3; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_1_bits_reg_idxw; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_wfd; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_fence; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_sfu; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_readmask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_writemask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_1_bits_wxd; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_1_bits_pc; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_ready; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_valid; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_2_bits_inst; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_wid; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_fp; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_branch; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_simt_stack; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_simt_stack_op; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_barrier; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_csr; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_reverse; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_sel_alu2; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_sel_alu1; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_isvec; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_sel_alu3; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_mask; // @[pipe.scala 54:27]
  wire [2:0] ibuffer2issue_io_in_2_bits_sel_imm; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_mem_unsigned; // @[pipe.scala 54:27]
  wire [5:0] ibuffer2issue_io_in_2_bits_alu_fn; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_mem; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_mem_cmd; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_2_bits_mop; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_2_bits_reg_idx1; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_2_bits_reg_idx2; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_2_bits_reg_idx3; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_2_bits_reg_idxw; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_wfd; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_fence; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_sfu; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_readmask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_writemask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_2_bits_wxd; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_2_bits_pc; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_ready; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_valid; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_3_bits_inst; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_wid; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_fp; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_branch; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_simt_stack; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_simt_stack_op; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_barrier; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_csr; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_reverse; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_sel_alu2; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_sel_alu1; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_isvec; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_sel_alu3; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_mask; // @[pipe.scala 54:27]
  wire [2:0] ibuffer2issue_io_in_3_bits_sel_imm; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_mem_unsigned; // @[pipe.scala 54:27]
  wire [5:0] ibuffer2issue_io_in_3_bits_alu_fn; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_mem; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_mem_cmd; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_in_3_bits_mop; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_3_bits_reg_idx1; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_3_bits_reg_idx2; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_3_bits_reg_idx3; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_in_3_bits_reg_idxw; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_wfd; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_fence; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_sfu; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_readmask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_writemask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_in_3_bits_wxd; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_in_3_bits_pc; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_ready; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_valid; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_out_bits_inst; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_wid; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_fp; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_branch; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_simt_stack; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_simt_stack_op; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_barrier; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_csr; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_reverse; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_sel_alu2; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_sel_alu1; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_isvec; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_sel_alu3; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_mask; // @[pipe.scala 54:27]
  wire [2:0] ibuffer2issue_io_out_bits_sel_imm; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_mem_unsigned; // @[pipe.scala 54:27]
  wire [5:0] ibuffer2issue_io_out_bits_alu_fn; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_mem; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_mem_cmd; // @[pipe.scala 54:27]
  wire [1:0] ibuffer2issue_io_out_bits_mop; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_out_bits_reg_idx1; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_out_bits_reg_idx2; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_out_bits_reg_idx3; // @[pipe.scala 54:27]
  wire [4:0] ibuffer2issue_io_out_bits_reg_idxw; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_wfd; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_fence; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_sfu; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_readmask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_writemask; // @[pipe.scala 54:27]
  wire  ibuffer2issue_io_out_bits_wxd; // @[pipe.scala 54:27]
  wire [31:0] ibuffer2issue_io_out_bits_pc; // @[pipe.scala 54:27]
  wire  exe_data_clock; // @[pipe.scala 55:22]
  wire  exe_data_reset; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_ready; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_valid; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_0; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_1; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_2; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_3; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_4; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_5; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_6; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in1_7; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_0; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_1; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_2; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_3; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_4; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_5; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_6; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in2_7; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_0; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_1; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_2; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_3; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_4; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_5; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_6; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_in3_7; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_0; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_1; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_2; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_3; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_4; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_5; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_6; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_mask_7; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_ctrl_inst; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_enq_bits_ctrl_wid; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_fp; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_enq_bits_ctrl_branch; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_simt_stack; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_simt_stack_op; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_barrier; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_enq_bits_ctrl_csr; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_reverse; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_isvec; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_mem_unsigned; // @[pipe.scala 55:22]
  wire [5:0] exe_data_io_enq_bits_ctrl_alu_fn; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_mem; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_enq_bits_ctrl_mem_cmd; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_enq_bits_ctrl_mop; // @[pipe.scala 55:22]
  wire [4:0] exe_data_io_enq_bits_ctrl_reg_idxw; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_wfd; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_fence; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_sfu; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_readmask; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_writemask; // @[pipe.scala 55:22]
  wire  exe_data_io_enq_bits_ctrl_wxd; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_enq_bits_ctrl_pc; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_ready; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_valid; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_0; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_1; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_2; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_3; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_4; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_5; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_6; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in1_7; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_0; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_1; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_2; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_3; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_4; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_5; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_6; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in2_7; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_0; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_1; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_2; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_3; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_4; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_5; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_6; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_in3_7; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_0; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_1; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_2; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_3; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_4; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_5; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_6; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_mask_7; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_ctrl_inst; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_deq_bits_ctrl_wid; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_fp; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_deq_bits_ctrl_branch; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_simt_stack; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_simt_stack_op; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_barrier; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_deq_bits_ctrl_csr; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_reverse; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_isvec; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_mem_unsigned; // @[pipe.scala 55:22]
  wire [5:0] exe_data_io_deq_bits_ctrl_alu_fn; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_mem; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_deq_bits_ctrl_mem_cmd; // @[pipe.scala 55:22]
  wire [1:0] exe_data_io_deq_bits_ctrl_mop; // @[pipe.scala 55:22]
  wire [4:0] exe_data_io_deq_bits_ctrl_reg_idxw; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_wfd; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_fence; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_sfu; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_readmask; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_writemask; // @[pipe.scala 55:22]
  wire  exe_data_io_deq_bits_ctrl_wxd; // @[pipe.scala 55:22]
  wire [31:0] exe_data_io_deq_bits_ctrl_pc; // @[pipe.scala 55:22]
  wire  simt_stack_clock; // @[pipe.scala 56:24]
  wire  simt_stack_reset; // @[pipe.scala 56:24]
  wire  simt_stack_io_branch_ctl_ready; // @[pipe.scala 56:24]
  wire  simt_stack_io_branch_ctl_valid; // @[pipe.scala 56:24]
  wire  simt_stack_io_branch_ctl_bits_opcode; // @[pipe.scala 56:24]
  wire [1:0] simt_stack_io_branch_ctl_bits_wid; // @[pipe.scala 56:24]
  wire [31:0] simt_stack_io_branch_ctl_bits_PC_branch; // @[pipe.scala 56:24]
  wire [7:0] simt_stack_io_branch_ctl_bits_mask_init; // @[pipe.scala 56:24]
  wire  simt_stack_io_if_mask_ready; // @[pipe.scala 56:24]
  wire  simt_stack_io_if_mask_valid; // @[pipe.scala 56:24]
  wire [7:0] simt_stack_io_if_mask_bits_if_mask; // @[pipe.scala 56:24]
  wire [1:0] simt_stack_io_if_mask_bits_wid; // @[pipe.scala 56:24]
  wire [1:0] simt_stack_io_input_wid; // @[pipe.scala 56:24]
  wire [7:0] simt_stack_io_out_mask; // @[pipe.scala 56:24]
  wire  simt_stack_io_complete_valid; // @[pipe.scala 56:24]
  wire [1:0] simt_stack_io_complete_bits; // @[pipe.scala 56:24]
  wire  simt_stack_io_fetch_ctl_ready; // @[pipe.scala 56:24]
  wire  simt_stack_io_fetch_ctl_valid; // @[pipe.scala 56:24]
  wire [1:0] simt_stack_io_fetch_ctl_bits_wid; // @[pipe.scala 56:24]
  wire  simt_stack_io_fetch_ctl_bits_jump; // @[pipe.scala 56:24]
  wire [31:0] simt_stack_io_fetch_ctl_bits_new_pc; // @[pipe.scala 56:24]
  wire  branch_back_io_out_ready; // @[pipe.scala 57:25]
  wire  branch_back_io_out_valid; // @[pipe.scala 57:25]
  wire [1:0] branch_back_io_out_bits_wid; // @[pipe.scala 57:25]
  wire  branch_back_io_out_bits_jump; // @[pipe.scala 57:25]
  wire [31:0] branch_back_io_out_bits_new_pc; // @[pipe.scala 57:25]
  wire  branch_back_io_in0_ready; // @[pipe.scala 57:25]
  wire  branch_back_io_in0_valid; // @[pipe.scala 57:25]
  wire [1:0] branch_back_io_in0_bits_wid; // @[pipe.scala 57:25]
  wire  branch_back_io_in0_bits_jump; // @[pipe.scala 57:25]
  wire [31:0] branch_back_io_in0_bits_new_pc; // @[pipe.scala 57:25]
  wire  branch_back_io_in1_ready; // @[pipe.scala 57:25]
  wire  branch_back_io_in1_valid; // @[pipe.scala 57:25]
  wire [1:0] branch_back_io_in1_bits_wid; // @[pipe.scala 57:25]
  wire  branch_back_io_in1_bits_jump; // @[pipe.scala 57:25]
  wire [31:0] branch_back_io_in1_bits_new_pc; // @[pipe.scala 57:25]
  wire  csrfile_clock; // @[pipe.scala 58:21]
  wire  csrfile_reset; // @[pipe.scala 58:21]
  wire  csrfile_io_in_ready; // @[pipe.scala 58:21]
  wire  csrfile_io_in_valid; // @[pipe.scala 58:21]
  wire [31:0] csrfile_io_in_bits_ctrl_inst; // @[pipe.scala 58:21]
  wire [1:0] csrfile_io_in_bits_ctrl_wid; // @[pipe.scala 58:21]
  wire [1:0] csrfile_io_in_bits_ctrl_csr; // @[pipe.scala 58:21]
  wire  csrfile_io_in_bits_ctrl_isvec; // @[pipe.scala 58:21]
  wire [4:0] csrfile_io_in_bits_ctrl_reg_idxw; // @[pipe.scala 58:21]
  wire  csrfile_io_in_bits_ctrl_wxd; // @[pipe.scala 58:21]
  wire [31:0] csrfile_io_in_bits_in1; // @[pipe.scala 58:21]
  wire  csrfile_io_out_ready; // @[pipe.scala 58:21]
  wire  csrfile_io_out_valid; // @[pipe.scala 58:21]
  wire [31:0] csrfile_io_out_bits_wb_wxd_rd; // @[pipe.scala 58:21]
  wire  csrfile_io_out_bits_wxd; // @[pipe.scala 58:21]
  wire [4:0] csrfile_io_out_bits_reg_idxw; // @[pipe.scala 58:21]
  wire [1:0] csrfile_io_out_bits_warp_id; // @[pipe.scala 58:21]
  wire [1:0] csrfile_io_frm_wid; // @[pipe.scala 58:21]
  wire [2:0] csrfile_io_frm; // @[pipe.scala 58:21]
  wire  csrfile_io_CTA2csr_valid; // @[pipe.scala 58:21]
  wire [2:0] csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[pipe.scala 58:21]
  wire [9:0] csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[pipe.scala 58:21]
  wire [12:0] csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[pipe.scala 58:21]
  wire [12:0] csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[pipe.scala 58:21]
  wire [4:0] csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[pipe.scala 58:21]
  wire [12:0] csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[pipe.scala 58:21]
  wire [1:0] csrfile_io_CTA2csr_bits_wid; // @[pipe.scala 58:21]
  wire  _warp_sche_io_issued_warp_valid_T = exe_data_io_enq_ready & exe_data_io_enq_valid; // @[Decoupled.scala 50:35]
  wire  scoreb_1_delay = Scoreboard_1_io_delay; // @[pipe.scala 52:{21,21}]
  wire  scoreb_0_delay = Scoreboard_io_delay; // @[pipe.scala 52:{21,21}]
  wire [1:0] warp_sche_io_scoreboard_busy_lo = {scoreb_1_delay,scoreb_0_delay}; // @[pipe.scala 77:70]
  wire  scoreb_3_delay = Scoreboard_3_io_delay; // @[pipe.scala 52:{21,21}]
  wire  scoreb_2_delay = Scoreboard_2_io_delay; // @[pipe.scala 52:{21,21}]
  wire [1:0] warp_sche_io_scoreboard_busy_hi = {scoreb_3_delay,scoreb_2_delay}; // @[pipe.scala 77:70]
  wire  _T_1 = control_io_control_alu_fn == 6'h3f & ibuffer_io_in_valid; // @[pipe.scala 101:41]
  wire  _T_3 = ~reset; // @[pipe.scala 102:11]
  wire  _ibuffer_ready_1_T_1 = ibuffer_io_out_1_bits_isvec & ibuffer_io_out_1_bits_simt_stack; // @[pipe.scala 129:27]
  wire  _ibuffer_ready_1_T_6 = ibuffer_io_out_1_bits_barrier ? warp_sche_io_warp_control_ready : alu_io_in_ready; // @[pipe.scala 132:22]
  wire  _ibuffer_ready_1_T_7 = ibuffer_io_out_1_bits_isvec ? valu_io_in_ready : _ibuffer_ready_1_T_6; // @[pipe.scala 131:20]
  wire  _ibuffer_ready_1_T_8 = _ibuffer_ready_1_T_1 ? simt_stack_io_branch_ctl_ready : _ibuffer_ready_1_T_7; // @[pipe.scala 130:18]
  wire  _ibuffer_ready_1_T_9 = ibuffer_io_out_1_bits_isvec & ibuffer_io_out_1_bits_simt_stack & ~
    ibuffer_io_out_1_bits_simt_stack_op ? valu_io_in_ready & simt_stack_io_branch_ctl_ready : _ibuffer_ready_1_T_8; // @[pipe.scala 129:16]
  wire  _ibuffer_ready_1_T_10 = ibuffer_io_out_1_bits_mem ? lsu_io_lsu_req_ready : _ibuffer_ready_1_T_9; // @[pipe.scala 128:14]
  wire  _ibuffer_ready_1_T_11 = |ibuffer_io_out_1_bits_csr ? csrfile_io_in_ready : _ibuffer_ready_1_T_10; // @[pipe.scala 127:12]
  wire  _ibuffer_ready_1_T_12 = ibuffer_io_out_1_bits_fp ? fpu_io_in_ready : _ibuffer_ready_1_T_11; // @[pipe.scala 126:10]
  wire  ibuffer_ready_1 = ibuffer_io_out_1_bits_sfu ? sfu_io_in_ready : _ibuffer_ready_1_T_12; // @[pipe.scala 125:26]
  wire  _ibuffer_ready_0_T_1 = ibuffer_io_out_0_bits_isvec & ibuffer_io_out_0_bits_simt_stack; // @[pipe.scala 129:27]
  wire  _ibuffer_ready_0_T_6 = ibuffer_io_out_0_bits_barrier ? warp_sche_io_warp_control_ready : alu_io_in_ready; // @[pipe.scala 132:22]
  wire  _ibuffer_ready_0_T_7 = ibuffer_io_out_0_bits_isvec ? valu_io_in_ready : _ibuffer_ready_0_T_6; // @[pipe.scala 131:20]
  wire  _ibuffer_ready_0_T_8 = _ibuffer_ready_0_T_1 ? simt_stack_io_branch_ctl_ready : _ibuffer_ready_0_T_7; // @[pipe.scala 130:18]
  wire  _ibuffer_ready_0_T_9 = ibuffer_io_out_0_bits_isvec & ibuffer_io_out_0_bits_simt_stack & ~
    ibuffer_io_out_0_bits_simt_stack_op ? valu_io_in_ready & simt_stack_io_branch_ctl_ready : _ibuffer_ready_0_T_8; // @[pipe.scala 129:16]
  wire  _ibuffer_ready_0_T_10 = ibuffer_io_out_0_bits_mem ? lsu_io_lsu_req_ready : _ibuffer_ready_0_T_9; // @[pipe.scala 128:14]
  wire  _ibuffer_ready_0_T_11 = |ibuffer_io_out_0_bits_csr ? csrfile_io_in_ready : _ibuffer_ready_0_T_10; // @[pipe.scala 127:12]
  wire  _ibuffer_ready_0_T_12 = ibuffer_io_out_0_bits_fp ? fpu_io_in_ready : _ibuffer_ready_0_T_11; // @[pipe.scala 126:10]
  wire  ibuffer_ready_0 = ibuffer_io_out_0_bits_sfu ? sfu_io_in_ready : _ibuffer_ready_0_T_12; // @[pipe.scala 125:26]
  wire  _ibuffer_ready_3_T_1 = ibuffer_io_out_3_bits_isvec & ibuffer_io_out_3_bits_simt_stack; // @[pipe.scala 129:27]
  wire  _ibuffer_ready_3_T_6 = ibuffer_io_out_3_bits_barrier ? warp_sche_io_warp_control_ready : alu_io_in_ready; // @[pipe.scala 132:22]
  wire  _ibuffer_ready_3_T_7 = ibuffer_io_out_3_bits_isvec ? valu_io_in_ready : _ibuffer_ready_3_T_6; // @[pipe.scala 131:20]
  wire  _ibuffer_ready_3_T_8 = _ibuffer_ready_3_T_1 ? simt_stack_io_branch_ctl_ready : _ibuffer_ready_3_T_7; // @[pipe.scala 130:18]
  wire  _ibuffer_ready_3_T_9 = ibuffer_io_out_3_bits_isvec & ibuffer_io_out_3_bits_simt_stack & ~
    ibuffer_io_out_3_bits_simt_stack_op ? valu_io_in_ready & simt_stack_io_branch_ctl_ready : _ibuffer_ready_3_T_8; // @[pipe.scala 129:16]
  wire  _ibuffer_ready_3_T_10 = ibuffer_io_out_3_bits_mem ? lsu_io_lsu_req_ready : _ibuffer_ready_3_T_9; // @[pipe.scala 128:14]
  wire  _ibuffer_ready_3_T_11 = |ibuffer_io_out_3_bits_csr ? csrfile_io_in_ready : _ibuffer_ready_3_T_10; // @[pipe.scala 127:12]
  wire  _ibuffer_ready_3_T_12 = ibuffer_io_out_3_bits_fp ? fpu_io_in_ready : _ibuffer_ready_3_T_11; // @[pipe.scala 126:10]
  wire  ibuffer_ready_3 = ibuffer_io_out_3_bits_sfu ? sfu_io_in_ready : _ibuffer_ready_3_T_12; // @[pipe.scala 125:26]
  wire  _ibuffer_ready_2_T_1 = ibuffer_io_out_2_bits_isvec & ibuffer_io_out_2_bits_simt_stack; // @[pipe.scala 129:27]
  wire  _ibuffer_ready_2_T_6 = ibuffer_io_out_2_bits_barrier ? warp_sche_io_warp_control_ready : alu_io_in_ready; // @[pipe.scala 132:22]
  wire  _ibuffer_ready_2_T_7 = ibuffer_io_out_2_bits_isvec ? valu_io_in_ready : _ibuffer_ready_2_T_6; // @[pipe.scala 131:20]
  wire  _ibuffer_ready_2_T_8 = _ibuffer_ready_2_T_1 ? simt_stack_io_branch_ctl_ready : _ibuffer_ready_2_T_7; // @[pipe.scala 130:18]
  wire  _ibuffer_ready_2_T_9 = ibuffer_io_out_2_bits_isvec & ibuffer_io_out_2_bits_simt_stack & ~
    ibuffer_io_out_2_bits_simt_stack_op ? valu_io_in_ready & simt_stack_io_branch_ctl_ready : _ibuffer_ready_2_T_8; // @[pipe.scala 129:16]
  wire  _ibuffer_ready_2_T_10 = ibuffer_io_out_2_bits_mem ? lsu_io_lsu_req_ready : _ibuffer_ready_2_T_9; // @[pipe.scala 128:14]
  wire  _ibuffer_ready_2_T_11 = |ibuffer_io_out_2_bits_csr ? csrfile_io_in_ready : _ibuffer_ready_2_T_10; // @[pipe.scala 127:12]
  wire  _ibuffer_ready_2_T_12 = ibuffer_io_out_2_bits_fp ? fpu_io_in_ready : _ibuffer_ready_2_T_11; // @[pipe.scala 126:10]
  wire  ibuffer_ready_2 = ibuffer_io_out_2_bits_sfu ? sfu_io_in_ready : _ibuffer_ready_2_T_12; // @[pipe.scala 125:26]
  wire [3:0] _warp_sche_io_exe_busy_T = {ibuffer_ready_3,ibuffer_ready_2,ibuffer_ready_1,ibuffer_ready_0}; // @[pipe.scala 116:48]
  wire  _T_4 = warp_sche_io_branch_ready & warp_sche_io_branch_valid; // @[Decoupled.scala 50:35]
  wire  _T_7 = warp_sche_io_warp_control_ready & warp_sche_io_warp_control_valid; // @[Decoupled.scala 50:35]
  wire  _T_11 = simt_stack_io_complete_valid & simt_stack_io_complete_bits == 2'h0; // @[pipe.scala 145:44]
  wire  _GEN_1 = _T_7 & warp_sche_io_warp_control_bits_ctrl_wid == 2'h0 | _T_11; // @[pipe.scala 144:{104,122}]
  wire  _T_19 = simt_stack_io_complete_valid & simt_stack_io_complete_bits == 2'h1; // @[pipe.scala 145:44]
  wire  _GEN_4 = _T_7 & warp_sche_io_warp_control_bits_ctrl_wid == 2'h1 | _T_19; // @[pipe.scala 144:{104,122}]
  wire  _T_27 = simt_stack_io_complete_valid & simt_stack_io_complete_bits == 2'h2; // @[pipe.scala 145:44]
  wire  _GEN_7 = _T_7 & warp_sche_io_warp_control_bits_ctrl_wid == 2'h2 | _T_27; // @[pipe.scala 144:{104,122}]
  wire  _T_35 = simt_stack_io_complete_valid & simt_stack_io_complete_bits == 2'h3; // @[pipe.scala 145:44]
  wire  _GEN_10 = _T_7 & warp_sche_io_warp_control_bits_ctrl_wid == 2'h3 | _T_35; // @[pipe.scala 144:{104,122}]
  wire  _scoreb_wb_x_fire_T = wb_io_out_x_ready & wb_io_out_x_valid; // @[Decoupled.scala 50:35]
  wire  _scoreb_wb_v_fire_T = wb_io_out_v_ready & wb_io_out_v_valid; // @[Decoupled.scala 50:35]
  wire  _T_42 = exe_data_io_deq_ready & exe_data_io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _T_53 = (exe_data_io_deq_bits_ctrl_wid == 2'h0 | exe_data_io_deq_bits_ctrl_wid == 2'h1) & _T_42 &
    exe_data_io_deq_bits_ctrl_alu_fn == 6'h6; // @[pipe.scala 186:115]
  warp_scheduler warp_sche ( // @[pipe.scala 39:23]
    .clock(warp_sche_clock),
    .reset(warp_sche_reset),
    .io_pc_reset(warp_sche_io_pc_reset),
    .io_warpReq_ready(warp_sche_io_warpReq_ready),
    .io_warpReq_valid(warp_sche_io_warpReq_valid),
    .io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count(warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch(warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch
      ),
    .io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch(warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch(
      warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch(
      warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch),
    .io_warpReq_bits_wid(warp_sche_io_warpReq_bits_wid),
    .io_warpRsp_valid(warp_sche_io_warpRsp_valid),
    .io_warpRsp_bits_wid(warp_sche_io_warpRsp_bits_wid),
    .io_wg_id_lookup(warp_sche_io_wg_id_lookup),
    .io_wg_id_tag(warp_sche_io_wg_id_tag),
    .io_pc_req_valid(warp_sche_io_pc_req_valid),
    .io_pc_req_bits_addr(warp_sche_io_pc_req_bits_addr),
    .io_pc_req_bits_warpid(warp_sche_io_pc_req_bits_warpid),
    .io_pc_rsp_valid(warp_sche_io_pc_rsp_valid),
    .io_pc_rsp_bits_addr(warp_sche_io_pc_rsp_bits_addr),
    .io_pc_rsp_bits_warpid(warp_sche_io_pc_rsp_bits_warpid),
    .io_pc_rsp_bits_status(warp_sche_io_pc_rsp_bits_status),
    .io_branch_ready(warp_sche_io_branch_ready),
    .io_branch_valid(warp_sche_io_branch_valid),
    .io_branch_bits_wid(warp_sche_io_branch_bits_wid),
    .io_branch_bits_jump(warp_sche_io_branch_bits_jump),
    .io_branch_bits_new_pc(warp_sche_io_branch_bits_new_pc),
    .io_warp_control_ready(warp_sche_io_warp_control_ready),
    .io_warp_control_valid(warp_sche_io_warp_control_valid),
    .io_warp_control_bits_ctrl_wid(warp_sche_io_warp_control_bits_ctrl_wid),
    .io_warp_control_bits_ctrl_simt_stack_op(warp_sche_io_warp_control_bits_ctrl_simt_stack_op),
    .io_warp_control_bits_ctrl_barrier(warp_sche_io_warp_control_bits_ctrl_barrier),
    .io_scoreboard_busy(warp_sche_io_scoreboard_busy),
    .io_exe_busy(warp_sche_io_exe_busy),
    .io_pc_ibuffer_ready_0(warp_sche_io_pc_ibuffer_ready_0),
    .io_pc_ibuffer_ready_1(warp_sche_io_pc_ibuffer_ready_1),
    .io_pc_ibuffer_ready_2(warp_sche_io_pc_ibuffer_ready_2),
    .io_pc_ibuffer_ready_3(warp_sche_io_pc_ibuffer_ready_3),
    .io_warp_ready(warp_sche_io_warp_ready),
    .io_flush_valid(warp_sche_io_flush_valid),
    .io_flush_bits(warp_sche_io_flush_bits),
    .io_flushCache_valid(warp_sche_io_flushCache_valid),
    .io_flushCache_bits(warp_sche_io_flushCache_bits),
    .io_CTA2csr_valid(warp_sche_io_CTA2csr_valid),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count(warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch(warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch
      ),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch(warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch(
      warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch),
    .io_CTA2csr_bits_wid(warp_sche_io_CTA2csr_bits_wid)
  );
  Control control ( // @[pipe.scala 41:21]
    .io_inst(control_io_inst),
    .io_pc(control_io_pc),
    .io_wid(control_io_wid),
    .io_control_inst(control_io_control_inst),
    .io_control_wid(control_io_control_wid),
    .io_control_fp(control_io_control_fp),
    .io_control_branch(control_io_control_branch),
    .io_control_simt_stack(control_io_control_simt_stack),
    .io_control_simt_stack_op(control_io_control_simt_stack_op),
    .io_control_barrier(control_io_control_barrier),
    .io_control_csr(control_io_control_csr),
    .io_control_reverse(control_io_control_reverse),
    .io_control_sel_alu2(control_io_control_sel_alu2),
    .io_control_sel_alu1(control_io_control_sel_alu1),
    .io_control_isvec(control_io_control_isvec),
    .io_control_sel_alu3(control_io_control_sel_alu3),
    .io_control_mask(control_io_control_mask),
    .io_control_sel_imm(control_io_control_sel_imm),
    .io_control_mem_unsigned(control_io_control_mem_unsigned),
    .io_control_alu_fn(control_io_control_alu_fn),
    .io_control_mem(control_io_control_mem),
    .io_control_mem_cmd(control_io_control_mem_cmd),
    .io_control_mop(control_io_control_mop),
    .io_control_reg_idx1(control_io_control_reg_idx1),
    .io_control_reg_idx2(control_io_control_reg_idx2),
    .io_control_reg_idx3(control_io_control_reg_idx3),
    .io_control_reg_idxw(control_io_control_reg_idxw),
    .io_control_wfd(control_io_control_wfd),
    .io_control_fence(control_io_control_fence),
    .io_control_sfu(control_io_control_sfu),
    .io_control_readmask(control_io_control_readmask),
    .io_control_writemask(control_io_control_writemask),
    .io_control_wxd(control_io_control_wxd),
    .io_control_pc(control_io_control_pc)
  );
  operandCollector operand_collector ( // @[pipe.scala 42:31]
    .clock(operand_collector_clock),
    .io_control_inst(operand_collector_io_control_inst),
    .io_control_wid(operand_collector_io_control_wid),
    .io_control_branch(operand_collector_io_control_branch),
    .io_control_sel_alu2(operand_collector_io_control_sel_alu2),
    .io_control_sel_alu1(operand_collector_io_control_sel_alu1),
    .io_control_isvec(operand_collector_io_control_isvec),
    .io_control_sel_alu3(operand_collector_io_control_sel_alu3),
    .io_control_mask(operand_collector_io_control_mask),
    .io_control_sel_imm(operand_collector_io_control_sel_imm),
    .io_control_reg_idx1(operand_collector_io_control_reg_idx1),
    .io_control_reg_idx2(operand_collector_io_control_reg_idx2),
    .io_control_reg_idx3(operand_collector_io_control_reg_idx3),
    .io_control_pc(operand_collector_io_control_pc),
    .io_alu_src1_0(operand_collector_io_alu_src1_0),
    .io_alu_src1_1(operand_collector_io_alu_src1_1),
    .io_alu_src1_2(operand_collector_io_alu_src1_2),
    .io_alu_src1_3(operand_collector_io_alu_src1_3),
    .io_alu_src1_4(operand_collector_io_alu_src1_4),
    .io_alu_src1_5(operand_collector_io_alu_src1_5),
    .io_alu_src1_6(operand_collector_io_alu_src1_6),
    .io_alu_src1_7(operand_collector_io_alu_src1_7),
    .io_alu_src2_0(operand_collector_io_alu_src2_0),
    .io_alu_src2_1(operand_collector_io_alu_src2_1),
    .io_alu_src2_2(operand_collector_io_alu_src2_2),
    .io_alu_src2_3(operand_collector_io_alu_src2_3),
    .io_alu_src2_4(operand_collector_io_alu_src2_4),
    .io_alu_src2_5(operand_collector_io_alu_src2_5),
    .io_alu_src2_6(operand_collector_io_alu_src2_6),
    .io_alu_src2_7(operand_collector_io_alu_src2_7),
    .io_alu_src3_0(operand_collector_io_alu_src3_0),
    .io_alu_src3_1(operand_collector_io_alu_src3_1),
    .io_alu_src3_2(operand_collector_io_alu_src3_2),
    .io_alu_src3_3(operand_collector_io_alu_src3_3),
    .io_alu_src3_4(operand_collector_io_alu_src3_4),
    .io_alu_src3_5(operand_collector_io_alu_src3_5),
    .io_alu_src3_6(operand_collector_io_alu_src3_6),
    .io_alu_src3_7(operand_collector_io_alu_src3_7),
    .io_mask_0(operand_collector_io_mask_0),
    .io_mask_1(operand_collector_io_mask_1),
    .io_mask_2(operand_collector_io_mask_2),
    .io_mask_3(operand_collector_io_mask_3),
    .io_mask_4(operand_collector_io_mask_4),
    .io_mask_5(operand_collector_io_mask_5),
    .io_mask_6(operand_collector_io_mask_6),
    .io_mask_7(operand_collector_io_mask_7),
    .io_writeScalarCtrl_valid(operand_collector_io_writeScalarCtrl_valid),
    .io_writeScalarCtrl_bits_wb_wxd_rd(operand_collector_io_writeScalarCtrl_bits_wb_wxd_rd),
    .io_writeScalarCtrl_bits_wxd(operand_collector_io_writeScalarCtrl_bits_wxd),
    .io_writeScalarCtrl_bits_reg_idxw(operand_collector_io_writeScalarCtrl_bits_reg_idxw),
    .io_writeScalarCtrl_bits_warp_id(operand_collector_io_writeScalarCtrl_bits_warp_id),
    .io_writeVecCtrl_valid(operand_collector_io_writeVecCtrl_valid),
    .io_writeVecCtrl_bits_wb_wfd_rd_0(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_0),
    .io_writeVecCtrl_bits_wb_wfd_rd_1(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_1),
    .io_writeVecCtrl_bits_wb_wfd_rd_2(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_2),
    .io_writeVecCtrl_bits_wb_wfd_rd_3(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_3),
    .io_writeVecCtrl_bits_wb_wfd_rd_4(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_4),
    .io_writeVecCtrl_bits_wb_wfd_rd_5(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_5),
    .io_writeVecCtrl_bits_wb_wfd_rd_6(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_6),
    .io_writeVecCtrl_bits_wb_wfd_rd_7(operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_7),
    .io_writeVecCtrl_bits_wfd_mask_0(operand_collector_io_writeVecCtrl_bits_wfd_mask_0),
    .io_writeVecCtrl_bits_wfd_mask_1(operand_collector_io_writeVecCtrl_bits_wfd_mask_1),
    .io_writeVecCtrl_bits_wfd_mask_2(operand_collector_io_writeVecCtrl_bits_wfd_mask_2),
    .io_writeVecCtrl_bits_wfd_mask_3(operand_collector_io_writeVecCtrl_bits_wfd_mask_3),
    .io_writeVecCtrl_bits_wfd_mask_4(operand_collector_io_writeVecCtrl_bits_wfd_mask_4),
    .io_writeVecCtrl_bits_wfd_mask_5(operand_collector_io_writeVecCtrl_bits_wfd_mask_5),
    .io_writeVecCtrl_bits_wfd_mask_6(operand_collector_io_writeVecCtrl_bits_wfd_mask_6),
    .io_writeVecCtrl_bits_wfd_mask_7(operand_collector_io_writeVecCtrl_bits_wfd_mask_7),
    .io_writeVecCtrl_bits_wfd(operand_collector_io_writeVecCtrl_bits_wfd),
    .io_writeVecCtrl_bits_reg_idxw(operand_collector_io_writeVecCtrl_bits_reg_idxw),
    .io_writeVecCtrl_bits_warp_id(operand_collector_io_writeVecCtrl_bits_warp_id)
  );
  Issue issue ( // @[pipe.scala 43:19]
    .io_in_ready(issue_io_in_ready),
    .io_in_valid(issue_io_in_valid),
    .io_in_bits_in1_0(issue_io_in_bits_in1_0),
    .io_in_bits_in1_1(issue_io_in_bits_in1_1),
    .io_in_bits_in1_2(issue_io_in_bits_in1_2),
    .io_in_bits_in1_3(issue_io_in_bits_in1_3),
    .io_in_bits_in1_4(issue_io_in_bits_in1_4),
    .io_in_bits_in1_5(issue_io_in_bits_in1_5),
    .io_in_bits_in1_6(issue_io_in_bits_in1_6),
    .io_in_bits_in1_7(issue_io_in_bits_in1_7),
    .io_in_bits_in2_0(issue_io_in_bits_in2_0),
    .io_in_bits_in2_1(issue_io_in_bits_in2_1),
    .io_in_bits_in2_2(issue_io_in_bits_in2_2),
    .io_in_bits_in2_3(issue_io_in_bits_in2_3),
    .io_in_bits_in2_4(issue_io_in_bits_in2_4),
    .io_in_bits_in2_5(issue_io_in_bits_in2_5),
    .io_in_bits_in2_6(issue_io_in_bits_in2_6),
    .io_in_bits_in2_7(issue_io_in_bits_in2_7),
    .io_in_bits_in3_0(issue_io_in_bits_in3_0),
    .io_in_bits_in3_1(issue_io_in_bits_in3_1),
    .io_in_bits_in3_2(issue_io_in_bits_in3_2),
    .io_in_bits_in3_3(issue_io_in_bits_in3_3),
    .io_in_bits_in3_4(issue_io_in_bits_in3_4),
    .io_in_bits_in3_5(issue_io_in_bits_in3_5),
    .io_in_bits_in3_6(issue_io_in_bits_in3_6),
    .io_in_bits_in3_7(issue_io_in_bits_in3_7),
    .io_in_bits_mask_0(issue_io_in_bits_mask_0),
    .io_in_bits_mask_1(issue_io_in_bits_mask_1),
    .io_in_bits_mask_2(issue_io_in_bits_mask_2),
    .io_in_bits_mask_3(issue_io_in_bits_mask_3),
    .io_in_bits_mask_4(issue_io_in_bits_mask_4),
    .io_in_bits_mask_5(issue_io_in_bits_mask_5),
    .io_in_bits_mask_6(issue_io_in_bits_mask_6),
    .io_in_bits_mask_7(issue_io_in_bits_mask_7),
    .io_in_bits_ctrl_inst(issue_io_in_bits_ctrl_inst),
    .io_in_bits_ctrl_wid(issue_io_in_bits_ctrl_wid),
    .io_in_bits_ctrl_fp(issue_io_in_bits_ctrl_fp),
    .io_in_bits_ctrl_branch(issue_io_in_bits_ctrl_branch),
    .io_in_bits_ctrl_simt_stack(issue_io_in_bits_ctrl_simt_stack),
    .io_in_bits_ctrl_simt_stack_op(issue_io_in_bits_ctrl_simt_stack_op),
    .io_in_bits_ctrl_barrier(issue_io_in_bits_ctrl_barrier),
    .io_in_bits_ctrl_csr(issue_io_in_bits_ctrl_csr),
    .io_in_bits_ctrl_reverse(issue_io_in_bits_ctrl_reverse),
    .io_in_bits_ctrl_isvec(issue_io_in_bits_ctrl_isvec),
    .io_in_bits_ctrl_mem_unsigned(issue_io_in_bits_ctrl_mem_unsigned),
    .io_in_bits_ctrl_alu_fn(issue_io_in_bits_ctrl_alu_fn),
    .io_in_bits_ctrl_mem(issue_io_in_bits_ctrl_mem),
    .io_in_bits_ctrl_mem_cmd(issue_io_in_bits_ctrl_mem_cmd),
    .io_in_bits_ctrl_mop(issue_io_in_bits_ctrl_mop),
    .io_in_bits_ctrl_reg_idxw(issue_io_in_bits_ctrl_reg_idxw),
    .io_in_bits_ctrl_wfd(issue_io_in_bits_ctrl_wfd),
    .io_in_bits_ctrl_fence(issue_io_in_bits_ctrl_fence),
    .io_in_bits_ctrl_sfu(issue_io_in_bits_ctrl_sfu),
    .io_in_bits_ctrl_readmask(issue_io_in_bits_ctrl_readmask),
    .io_in_bits_ctrl_writemask(issue_io_in_bits_ctrl_writemask),
    .io_in_bits_ctrl_wxd(issue_io_in_bits_ctrl_wxd),
    .io_in_bits_ctrl_pc(issue_io_in_bits_ctrl_pc),
    .io_out_sALU_ready(issue_io_out_sALU_ready),
    .io_out_sALU_valid(issue_io_out_sALU_valid),
    .io_out_sALU_bits_in1(issue_io_out_sALU_bits_in1),
    .io_out_sALU_bits_in2(issue_io_out_sALU_bits_in2),
    .io_out_sALU_bits_in3(issue_io_out_sALU_bits_in3),
    .io_out_sALU_bits_ctrl_wid(issue_io_out_sALU_bits_ctrl_wid),
    .io_out_sALU_bits_ctrl_branch(issue_io_out_sALU_bits_ctrl_branch),
    .io_out_sALU_bits_ctrl_alu_fn(issue_io_out_sALU_bits_ctrl_alu_fn),
    .io_out_sALU_bits_ctrl_reg_idxw(issue_io_out_sALU_bits_ctrl_reg_idxw),
    .io_out_sALU_bits_ctrl_wxd(issue_io_out_sALU_bits_ctrl_wxd),
    .io_out_vALU_ready(issue_io_out_vALU_ready),
    .io_out_vALU_valid(issue_io_out_vALU_valid),
    .io_out_vALU_bits_in1_0(issue_io_out_vALU_bits_in1_0),
    .io_out_vALU_bits_in1_1(issue_io_out_vALU_bits_in1_1),
    .io_out_vALU_bits_in1_2(issue_io_out_vALU_bits_in1_2),
    .io_out_vALU_bits_in1_3(issue_io_out_vALU_bits_in1_3),
    .io_out_vALU_bits_in1_4(issue_io_out_vALU_bits_in1_4),
    .io_out_vALU_bits_in1_5(issue_io_out_vALU_bits_in1_5),
    .io_out_vALU_bits_in1_6(issue_io_out_vALU_bits_in1_6),
    .io_out_vALU_bits_in1_7(issue_io_out_vALU_bits_in1_7),
    .io_out_vALU_bits_in2_0(issue_io_out_vALU_bits_in2_0),
    .io_out_vALU_bits_in2_1(issue_io_out_vALU_bits_in2_1),
    .io_out_vALU_bits_in2_2(issue_io_out_vALU_bits_in2_2),
    .io_out_vALU_bits_in2_3(issue_io_out_vALU_bits_in2_3),
    .io_out_vALU_bits_in2_4(issue_io_out_vALU_bits_in2_4),
    .io_out_vALU_bits_in2_5(issue_io_out_vALU_bits_in2_5),
    .io_out_vALU_bits_in2_6(issue_io_out_vALU_bits_in2_6),
    .io_out_vALU_bits_in2_7(issue_io_out_vALU_bits_in2_7),
    .io_out_vALU_bits_in3_0(issue_io_out_vALU_bits_in3_0),
    .io_out_vALU_bits_in3_1(issue_io_out_vALU_bits_in3_1),
    .io_out_vALU_bits_in3_2(issue_io_out_vALU_bits_in3_2),
    .io_out_vALU_bits_in3_3(issue_io_out_vALU_bits_in3_3),
    .io_out_vALU_bits_in3_4(issue_io_out_vALU_bits_in3_4),
    .io_out_vALU_bits_in3_5(issue_io_out_vALU_bits_in3_5),
    .io_out_vALU_bits_in3_6(issue_io_out_vALU_bits_in3_6),
    .io_out_vALU_bits_in3_7(issue_io_out_vALU_bits_in3_7),
    .io_out_vALU_bits_mask_0(issue_io_out_vALU_bits_mask_0),
    .io_out_vALU_bits_mask_1(issue_io_out_vALU_bits_mask_1),
    .io_out_vALU_bits_mask_2(issue_io_out_vALU_bits_mask_2),
    .io_out_vALU_bits_mask_3(issue_io_out_vALU_bits_mask_3),
    .io_out_vALU_bits_mask_4(issue_io_out_vALU_bits_mask_4),
    .io_out_vALU_bits_mask_5(issue_io_out_vALU_bits_mask_5),
    .io_out_vALU_bits_mask_6(issue_io_out_vALU_bits_mask_6),
    .io_out_vALU_bits_mask_7(issue_io_out_vALU_bits_mask_7),
    .io_out_vALU_bits_ctrl_wid(issue_io_out_vALU_bits_ctrl_wid),
    .io_out_vALU_bits_ctrl_simt_stack(issue_io_out_vALU_bits_ctrl_simt_stack),
    .io_out_vALU_bits_ctrl_reverse(issue_io_out_vALU_bits_ctrl_reverse),
    .io_out_vALU_bits_ctrl_alu_fn(issue_io_out_vALU_bits_ctrl_alu_fn),
    .io_out_vALU_bits_ctrl_reg_idxw(issue_io_out_vALU_bits_ctrl_reg_idxw),
    .io_out_vALU_bits_ctrl_wfd(issue_io_out_vALU_bits_ctrl_wfd),
    .io_out_vALU_bits_ctrl_readmask(issue_io_out_vALU_bits_ctrl_readmask),
    .io_out_vALU_bits_ctrl_writemask(issue_io_out_vALU_bits_ctrl_writemask),
    .io_out_vFPU_ready(issue_io_out_vFPU_ready),
    .io_out_vFPU_valid(issue_io_out_vFPU_valid),
    .io_out_vFPU_bits_in1_0(issue_io_out_vFPU_bits_in1_0),
    .io_out_vFPU_bits_in1_1(issue_io_out_vFPU_bits_in1_1),
    .io_out_vFPU_bits_in1_2(issue_io_out_vFPU_bits_in1_2),
    .io_out_vFPU_bits_in1_3(issue_io_out_vFPU_bits_in1_3),
    .io_out_vFPU_bits_in1_4(issue_io_out_vFPU_bits_in1_4),
    .io_out_vFPU_bits_in1_5(issue_io_out_vFPU_bits_in1_5),
    .io_out_vFPU_bits_in1_6(issue_io_out_vFPU_bits_in1_6),
    .io_out_vFPU_bits_in1_7(issue_io_out_vFPU_bits_in1_7),
    .io_out_vFPU_bits_in2_0(issue_io_out_vFPU_bits_in2_0),
    .io_out_vFPU_bits_in2_1(issue_io_out_vFPU_bits_in2_1),
    .io_out_vFPU_bits_in2_2(issue_io_out_vFPU_bits_in2_2),
    .io_out_vFPU_bits_in2_3(issue_io_out_vFPU_bits_in2_3),
    .io_out_vFPU_bits_in2_4(issue_io_out_vFPU_bits_in2_4),
    .io_out_vFPU_bits_in2_5(issue_io_out_vFPU_bits_in2_5),
    .io_out_vFPU_bits_in2_6(issue_io_out_vFPU_bits_in2_6),
    .io_out_vFPU_bits_in2_7(issue_io_out_vFPU_bits_in2_7),
    .io_out_vFPU_bits_in3_0(issue_io_out_vFPU_bits_in3_0),
    .io_out_vFPU_bits_in3_1(issue_io_out_vFPU_bits_in3_1),
    .io_out_vFPU_bits_in3_2(issue_io_out_vFPU_bits_in3_2),
    .io_out_vFPU_bits_in3_3(issue_io_out_vFPU_bits_in3_3),
    .io_out_vFPU_bits_in3_4(issue_io_out_vFPU_bits_in3_4),
    .io_out_vFPU_bits_in3_5(issue_io_out_vFPU_bits_in3_5),
    .io_out_vFPU_bits_in3_6(issue_io_out_vFPU_bits_in3_6),
    .io_out_vFPU_bits_in3_7(issue_io_out_vFPU_bits_in3_7),
    .io_out_vFPU_bits_mask_0(issue_io_out_vFPU_bits_mask_0),
    .io_out_vFPU_bits_mask_1(issue_io_out_vFPU_bits_mask_1),
    .io_out_vFPU_bits_mask_2(issue_io_out_vFPU_bits_mask_2),
    .io_out_vFPU_bits_mask_3(issue_io_out_vFPU_bits_mask_3),
    .io_out_vFPU_bits_mask_4(issue_io_out_vFPU_bits_mask_4),
    .io_out_vFPU_bits_mask_5(issue_io_out_vFPU_bits_mask_5),
    .io_out_vFPU_bits_mask_6(issue_io_out_vFPU_bits_mask_6),
    .io_out_vFPU_bits_mask_7(issue_io_out_vFPU_bits_mask_7),
    .io_out_vFPU_bits_ctrl_wid(issue_io_out_vFPU_bits_ctrl_wid),
    .io_out_vFPU_bits_ctrl_reverse(issue_io_out_vFPU_bits_ctrl_reverse),
    .io_out_vFPU_bits_ctrl_alu_fn(issue_io_out_vFPU_bits_ctrl_alu_fn),
    .io_out_vFPU_bits_ctrl_reg_idxw(issue_io_out_vFPU_bits_ctrl_reg_idxw),
    .io_out_vFPU_bits_ctrl_wfd(issue_io_out_vFPU_bits_ctrl_wfd),
    .io_out_vFPU_bits_ctrl_wxd(issue_io_out_vFPU_bits_ctrl_wxd),
    .io_out_LSU_ready(issue_io_out_LSU_ready),
    .io_out_LSU_valid(issue_io_out_LSU_valid),
    .io_out_LSU_bits_in1_0(issue_io_out_LSU_bits_in1_0),
    .io_out_LSU_bits_in1_1(issue_io_out_LSU_bits_in1_1),
    .io_out_LSU_bits_in1_2(issue_io_out_LSU_bits_in1_2),
    .io_out_LSU_bits_in1_3(issue_io_out_LSU_bits_in1_3),
    .io_out_LSU_bits_in1_4(issue_io_out_LSU_bits_in1_4),
    .io_out_LSU_bits_in1_5(issue_io_out_LSU_bits_in1_5),
    .io_out_LSU_bits_in1_6(issue_io_out_LSU_bits_in1_6),
    .io_out_LSU_bits_in1_7(issue_io_out_LSU_bits_in1_7),
    .io_out_LSU_bits_in2_0(issue_io_out_LSU_bits_in2_0),
    .io_out_LSU_bits_in2_1(issue_io_out_LSU_bits_in2_1),
    .io_out_LSU_bits_in2_2(issue_io_out_LSU_bits_in2_2),
    .io_out_LSU_bits_in2_3(issue_io_out_LSU_bits_in2_3),
    .io_out_LSU_bits_in2_4(issue_io_out_LSU_bits_in2_4),
    .io_out_LSU_bits_in2_5(issue_io_out_LSU_bits_in2_5),
    .io_out_LSU_bits_in2_6(issue_io_out_LSU_bits_in2_6),
    .io_out_LSU_bits_in2_7(issue_io_out_LSU_bits_in2_7),
    .io_out_LSU_bits_in3_0(issue_io_out_LSU_bits_in3_0),
    .io_out_LSU_bits_in3_1(issue_io_out_LSU_bits_in3_1),
    .io_out_LSU_bits_in3_2(issue_io_out_LSU_bits_in3_2),
    .io_out_LSU_bits_in3_3(issue_io_out_LSU_bits_in3_3),
    .io_out_LSU_bits_in3_4(issue_io_out_LSU_bits_in3_4),
    .io_out_LSU_bits_in3_5(issue_io_out_LSU_bits_in3_5),
    .io_out_LSU_bits_in3_6(issue_io_out_LSU_bits_in3_6),
    .io_out_LSU_bits_in3_7(issue_io_out_LSU_bits_in3_7),
    .io_out_LSU_bits_mask_0(issue_io_out_LSU_bits_mask_0),
    .io_out_LSU_bits_mask_1(issue_io_out_LSU_bits_mask_1),
    .io_out_LSU_bits_mask_2(issue_io_out_LSU_bits_mask_2),
    .io_out_LSU_bits_mask_3(issue_io_out_LSU_bits_mask_3),
    .io_out_LSU_bits_mask_4(issue_io_out_LSU_bits_mask_4),
    .io_out_LSU_bits_mask_5(issue_io_out_LSU_bits_mask_5),
    .io_out_LSU_bits_mask_6(issue_io_out_LSU_bits_mask_6),
    .io_out_LSU_bits_mask_7(issue_io_out_LSU_bits_mask_7),
    .io_out_LSU_bits_ctrl_inst(issue_io_out_LSU_bits_ctrl_inst),
    .io_out_LSU_bits_ctrl_wid(issue_io_out_LSU_bits_ctrl_wid),
    .io_out_LSU_bits_ctrl_fp(issue_io_out_LSU_bits_ctrl_fp),
    .io_out_LSU_bits_ctrl_branch(issue_io_out_LSU_bits_ctrl_branch),
    .io_out_LSU_bits_ctrl_simt_stack(issue_io_out_LSU_bits_ctrl_simt_stack),
    .io_out_LSU_bits_ctrl_simt_stack_op(issue_io_out_LSU_bits_ctrl_simt_stack_op),
    .io_out_LSU_bits_ctrl_barrier(issue_io_out_LSU_bits_ctrl_barrier),
    .io_out_LSU_bits_ctrl_csr(issue_io_out_LSU_bits_ctrl_csr),
    .io_out_LSU_bits_ctrl_reverse(issue_io_out_LSU_bits_ctrl_reverse),
    .io_out_LSU_bits_ctrl_isvec(issue_io_out_LSU_bits_ctrl_isvec),
    .io_out_LSU_bits_ctrl_mem_unsigned(issue_io_out_LSU_bits_ctrl_mem_unsigned),
    .io_out_LSU_bits_ctrl_alu_fn(issue_io_out_LSU_bits_ctrl_alu_fn),
    .io_out_LSU_bits_ctrl_mem(issue_io_out_LSU_bits_ctrl_mem),
    .io_out_LSU_bits_ctrl_mem_cmd(issue_io_out_LSU_bits_ctrl_mem_cmd),
    .io_out_LSU_bits_ctrl_mop(issue_io_out_LSU_bits_ctrl_mop),
    .io_out_LSU_bits_ctrl_reg_idxw(issue_io_out_LSU_bits_ctrl_reg_idxw),
    .io_out_LSU_bits_ctrl_wfd(issue_io_out_LSU_bits_ctrl_wfd),
    .io_out_LSU_bits_ctrl_fence(issue_io_out_LSU_bits_ctrl_fence),
    .io_out_LSU_bits_ctrl_sfu(issue_io_out_LSU_bits_ctrl_sfu),
    .io_out_LSU_bits_ctrl_readmask(issue_io_out_LSU_bits_ctrl_readmask),
    .io_out_LSU_bits_ctrl_writemask(issue_io_out_LSU_bits_ctrl_writemask),
    .io_out_LSU_bits_ctrl_wxd(issue_io_out_LSU_bits_ctrl_wxd),
    .io_out_LSU_bits_ctrl_pc(issue_io_out_LSU_bits_ctrl_pc),
    .io_out_SFU_ready(issue_io_out_SFU_ready),
    .io_out_SFU_valid(issue_io_out_SFU_valid),
    .io_out_SFU_bits_in1_0(issue_io_out_SFU_bits_in1_0),
    .io_out_SFU_bits_in1_1(issue_io_out_SFU_bits_in1_1),
    .io_out_SFU_bits_in1_2(issue_io_out_SFU_bits_in1_2),
    .io_out_SFU_bits_in1_3(issue_io_out_SFU_bits_in1_3),
    .io_out_SFU_bits_in1_4(issue_io_out_SFU_bits_in1_4),
    .io_out_SFU_bits_in1_5(issue_io_out_SFU_bits_in1_5),
    .io_out_SFU_bits_in1_6(issue_io_out_SFU_bits_in1_6),
    .io_out_SFU_bits_in1_7(issue_io_out_SFU_bits_in1_7),
    .io_out_SFU_bits_in2_0(issue_io_out_SFU_bits_in2_0),
    .io_out_SFU_bits_in2_1(issue_io_out_SFU_bits_in2_1),
    .io_out_SFU_bits_in2_2(issue_io_out_SFU_bits_in2_2),
    .io_out_SFU_bits_in2_3(issue_io_out_SFU_bits_in2_3),
    .io_out_SFU_bits_in2_4(issue_io_out_SFU_bits_in2_4),
    .io_out_SFU_bits_in2_5(issue_io_out_SFU_bits_in2_5),
    .io_out_SFU_bits_in2_6(issue_io_out_SFU_bits_in2_6),
    .io_out_SFU_bits_in2_7(issue_io_out_SFU_bits_in2_7),
    .io_out_SFU_bits_mask_0(issue_io_out_SFU_bits_mask_0),
    .io_out_SFU_bits_mask_1(issue_io_out_SFU_bits_mask_1),
    .io_out_SFU_bits_mask_2(issue_io_out_SFU_bits_mask_2),
    .io_out_SFU_bits_mask_3(issue_io_out_SFU_bits_mask_3),
    .io_out_SFU_bits_mask_4(issue_io_out_SFU_bits_mask_4),
    .io_out_SFU_bits_mask_5(issue_io_out_SFU_bits_mask_5),
    .io_out_SFU_bits_mask_6(issue_io_out_SFU_bits_mask_6),
    .io_out_SFU_bits_mask_7(issue_io_out_SFU_bits_mask_7),
    .io_out_SFU_bits_ctrl_wid(issue_io_out_SFU_bits_ctrl_wid),
    .io_out_SFU_bits_ctrl_fp(issue_io_out_SFU_bits_ctrl_fp),
    .io_out_SFU_bits_ctrl_reverse(issue_io_out_SFU_bits_ctrl_reverse),
    .io_out_SFU_bits_ctrl_isvec(issue_io_out_SFU_bits_ctrl_isvec),
    .io_out_SFU_bits_ctrl_alu_fn(issue_io_out_SFU_bits_ctrl_alu_fn),
    .io_out_SFU_bits_ctrl_reg_idxw(issue_io_out_SFU_bits_ctrl_reg_idxw),
    .io_out_SFU_bits_ctrl_wfd(issue_io_out_SFU_bits_ctrl_wfd),
    .io_out_SFU_bits_ctrl_wxd(issue_io_out_SFU_bits_ctrl_wxd),
    .io_out_SIMT_ready(issue_io_out_SIMT_ready),
    .io_out_SIMT_valid(issue_io_out_SIMT_valid),
    .io_out_SIMT_bits_opcode(issue_io_out_SIMT_bits_opcode),
    .io_out_SIMT_bits_wid(issue_io_out_SIMT_bits_wid),
    .io_out_SIMT_bits_PC_branch(issue_io_out_SIMT_bits_PC_branch),
    .io_out_SIMT_bits_mask_init(issue_io_out_SIMT_bits_mask_init),
    .io_out_warpscheduler_ready(issue_io_out_warpscheduler_ready),
    .io_out_warpscheduler_valid(issue_io_out_warpscheduler_valid),
    .io_out_warpscheduler_bits_ctrl_wid(issue_io_out_warpscheduler_bits_ctrl_wid),
    .io_out_warpscheduler_bits_ctrl_simt_stack_op(issue_io_out_warpscheduler_bits_ctrl_simt_stack_op),
    .io_out_warpscheduler_bits_ctrl_barrier(issue_io_out_warpscheduler_bits_ctrl_barrier),
    .io_out_CSR_ready(issue_io_out_CSR_ready),
    .io_out_CSR_valid(issue_io_out_CSR_valid),
    .io_out_CSR_bits_ctrl_inst(issue_io_out_CSR_bits_ctrl_inst),
    .io_out_CSR_bits_ctrl_wid(issue_io_out_CSR_bits_ctrl_wid),
    .io_out_CSR_bits_ctrl_csr(issue_io_out_CSR_bits_ctrl_csr),
    .io_out_CSR_bits_ctrl_isvec(issue_io_out_CSR_bits_ctrl_isvec),
    .io_out_CSR_bits_ctrl_reg_idxw(issue_io_out_CSR_bits_ctrl_reg_idxw),
    .io_out_CSR_bits_ctrl_wxd(issue_io_out_CSR_bits_ctrl_wxd),
    .io_out_CSR_bits_in1(issue_io_out_CSR_bits_in1)
  );
  ALUexe alu ( // @[pipe.scala 44:17]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_ready(alu_io_in_ready),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_in1(alu_io_in_bits_in1),
    .io_in_bits_in2(alu_io_in_bits_in2),
    .io_in_bits_in3(alu_io_in_bits_in3),
    .io_in_bits_ctrl_wid(alu_io_in_bits_ctrl_wid),
    .io_in_bits_ctrl_branch(alu_io_in_bits_ctrl_branch),
    .io_in_bits_ctrl_alu_fn(alu_io_in_bits_ctrl_alu_fn),
    .io_in_bits_ctrl_reg_idxw(alu_io_in_bits_ctrl_reg_idxw),
    .io_in_bits_ctrl_wxd(alu_io_in_bits_ctrl_wxd),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits_wb_wxd_rd(alu_io_out_bits_wb_wxd_rd),
    .io_out_bits_wxd(alu_io_out_bits_wxd),
    .io_out_bits_reg_idxw(alu_io_out_bits_reg_idxw),
    .io_out_bits_warp_id(alu_io_out_bits_warp_id),
    .io_out2br_ready(alu_io_out2br_ready),
    .io_out2br_valid(alu_io_out2br_valid),
    .io_out2br_bits_wid(alu_io_out2br_bits_wid),
    .io_out2br_bits_jump(alu_io_out2br_bits_jump),
    .io_out2br_bits_new_pc(alu_io_out2br_bits_new_pc)
  );
  vALUexe valu ( // @[pipe.scala 45:18]
    .clock(valu_clock),
    .reset(valu_reset),
    .io_in_ready(valu_io_in_ready),
    .io_in_valid(valu_io_in_valid),
    .io_in_bits_in1_0(valu_io_in_bits_in1_0),
    .io_in_bits_in1_1(valu_io_in_bits_in1_1),
    .io_in_bits_in1_2(valu_io_in_bits_in1_2),
    .io_in_bits_in1_3(valu_io_in_bits_in1_3),
    .io_in_bits_in1_4(valu_io_in_bits_in1_4),
    .io_in_bits_in1_5(valu_io_in_bits_in1_5),
    .io_in_bits_in1_6(valu_io_in_bits_in1_6),
    .io_in_bits_in1_7(valu_io_in_bits_in1_7),
    .io_in_bits_in2_0(valu_io_in_bits_in2_0),
    .io_in_bits_in2_1(valu_io_in_bits_in2_1),
    .io_in_bits_in2_2(valu_io_in_bits_in2_2),
    .io_in_bits_in2_3(valu_io_in_bits_in2_3),
    .io_in_bits_in2_4(valu_io_in_bits_in2_4),
    .io_in_bits_in2_5(valu_io_in_bits_in2_5),
    .io_in_bits_in2_6(valu_io_in_bits_in2_6),
    .io_in_bits_in2_7(valu_io_in_bits_in2_7),
    .io_in_bits_in3_0(valu_io_in_bits_in3_0),
    .io_in_bits_in3_1(valu_io_in_bits_in3_1),
    .io_in_bits_in3_2(valu_io_in_bits_in3_2),
    .io_in_bits_in3_3(valu_io_in_bits_in3_3),
    .io_in_bits_in3_4(valu_io_in_bits_in3_4),
    .io_in_bits_in3_5(valu_io_in_bits_in3_5),
    .io_in_bits_in3_6(valu_io_in_bits_in3_6),
    .io_in_bits_in3_7(valu_io_in_bits_in3_7),
    .io_in_bits_mask_0(valu_io_in_bits_mask_0),
    .io_in_bits_mask_1(valu_io_in_bits_mask_1),
    .io_in_bits_mask_2(valu_io_in_bits_mask_2),
    .io_in_bits_mask_3(valu_io_in_bits_mask_3),
    .io_in_bits_mask_4(valu_io_in_bits_mask_4),
    .io_in_bits_mask_5(valu_io_in_bits_mask_5),
    .io_in_bits_mask_6(valu_io_in_bits_mask_6),
    .io_in_bits_mask_7(valu_io_in_bits_mask_7),
    .io_in_bits_ctrl_wid(valu_io_in_bits_ctrl_wid),
    .io_in_bits_ctrl_simt_stack(valu_io_in_bits_ctrl_simt_stack),
    .io_in_bits_ctrl_reverse(valu_io_in_bits_ctrl_reverse),
    .io_in_bits_ctrl_alu_fn(valu_io_in_bits_ctrl_alu_fn),
    .io_in_bits_ctrl_reg_idxw(valu_io_in_bits_ctrl_reg_idxw),
    .io_in_bits_ctrl_wfd(valu_io_in_bits_ctrl_wfd),
    .io_in_bits_ctrl_readmask(valu_io_in_bits_ctrl_readmask),
    .io_in_bits_ctrl_writemask(valu_io_in_bits_ctrl_writemask),
    .io_out_valid(valu_io_out_valid),
    .io_out_bits_wb_wfd_rd_0(valu_io_out_bits_wb_wfd_rd_0),
    .io_out_bits_wb_wfd_rd_1(valu_io_out_bits_wb_wfd_rd_1),
    .io_out_bits_wb_wfd_rd_2(valu_io_out_bits_wb_wfd_rd_2),
    .io_out_bits_wb_wfd_rd_3(valu_io_out_bits_wb_wfd_rd_3),
    .io_out_bits_wb_wfd_rd_4(valu_io_out_bits_wb_wfd_rd_4),
    .io_out_bits_wb_wfd_rd_5(valu_io_out_bits_wb_wfd_rd_5),
    .io_out_bits_wb_wfd_rd_6(valu_io_out_bits_wb_wfd_rd_6),
    .io_out_bits_wb_wfd_rd_7(valu_io_out_bits_wb_wfd_rd_7),
    .io_out_bits_wfd_mask_0(valu_io_out_bits_wfd_mask_0),
    .io_out_bits_wfd_mask_1(valu_io_out_bits_wfd_mask_1),
    .io_out_bits_wfd_mask_2(valu_io_out_bits_wfd_mask_2),
    .io_out_bits_wfd_mask_3(valu_io_out_bits_wfd_mask_3),
    .io_out_bits_wfd_mask_4(valu_io_out_bits_wfd_mask_4),
    .io_out_bits_wfd_mask_5(valu_io_out_bits_wfd_mask_5),
    .io_out_bits_wfd_mask_6(valu_io_out_bits_wfd_mask_6),
    .io_out_bits_wfd_mask_7(valu_io_out_bits_wfd_mask_7),
    .io_out_bits_wfd(valu_io_out_bits_wfd),
    .io_out_bits_reg_idxw(valu_io_out_bits_reg_idxw),
    .io_out_bits_warp_id(valu_io_out_bits_warp_id),
    .io_out2simt_stack_ready(valu_io_out2simt_stack_ready),
    .io_out2simt_stack_valid(valu_io_out2simt_stack_valid),
    .io_out2simt_stack_bits_if_mask(valu_io_out2simt_stack_bits_if_mask),
    .io_out2simt_stack_bits_wid(valu_io_out2simt_stack_bits_wid)
  );
  FPUexe fpu ( // @[pipe.scala 46:17]
    .clock(fpu_clock),
    .reset(fpu_reset),
    .io_in_ready(fpu_io_in_ready),
    .io_in_valid(fpu_io_in_valid),
    .io_in_bits_in1_0(fpu_io_in_bits_in1_0),
    .io_in_bits_in1_1(fpu_io_in_bits_in1_1),
    .io_in_bits_in1_2(fpu_io_in_bits_in1_2),
    .io_in_bits_in1_3(fpu_io_in_bits_in1_3),
    .io_in_bits_in1_4(fpu_io_in_bits_in1_4),
    .io_in_bits_in1_5(fpu_io_in_bits_in1_5),
    .io_in_bits_in1_6(fpu_io_in_bits_in1_6),
    .io_in_bits_in1_7(fpu_io_in_bits_in1_7),
    .io_in_bits_in2_0(fpu_io_in_bits_in2_0),
    .io_in_bits_in2_1(fpu_io_in_bits_in2_1),
    .io_in_bits_in2_2(fpu_io_in_bits_in2_2),
    .io_in_bits_in2_3(fpu_io_in_bits_in2_3),
    .io_in_bits_in2_4(fpu_io_in_bits_in2_4),
    .io_in_bits_in2_5(fpu_io_in_bits_in2_5),
    .io_in_bits_in2_6(fpu_io_in_bits_in2_6),
    .io_in_bits_in2_7(fpu_io_in_bits_in2_7),
    .io_in_bits_in3_0(fpu_io_in_bits_in3_0),
    .io_in_bits_in3_1(fpu_io_in_bits_in3_1),
    .io_in_bits_in3_2(fpu_io_in_bits_in3_2),
    .io_in_bits_in3_3(fpu_io_in_bits_in3_3),
    .io_in_bits_in3_4(fpu_io_in_bits_in3_4),
    .io_in_bits_in3_5(fpu_io_in_bits_in3_5),
    .io_in_bits_in3_6(fpu_io_in_bits_in3_6),
    .io_in_bits_in3_7(fpu_io_in_bits_in3_7),
    .io_in_bits_mask_0(fpu_io_in_bits_mask_0),
    .io_in_bits_mask_1(fpu_io_in_bits_mask_1),
    .io_in_bits_mask_2(fpu_io_in_bits_mask_2),
    .io_in_bits_mask_3(fpu_io_in_bits_mask_3),
    .io_in_bits_mask_4(fpu_io_in_bits_mask_4),
    .io_in_bits_mask_5(fpu_io_in_bits_mask_5),
    .io_in_bits_mask_6(fpu_io_in_bits_mask_6),
    .io_in_bits_mask_7(fpu_io_in_bits_mask_7),
    .io_in_bits_ctrl_wid(fpu_io_in_bits_ctrl_wid),
    .io_in_bits_ctrl_reverse(fpu_io_in_bits_ctrl_reverse),
    .io_in_bits_ctrl_alu_fn(fpu_io_in_bits_ctrl_alu_fn),
    .io_in_bits_ctrl_reg_idxw(fpu_io_in_bits_ctrl_reg_idxw),
    .io_in_bits_ctrl_wfd(fpu_io_in_bits_ctrl_wfd),
    .io_in_bits_ctrl_wxd(fpu_io_in_bits_ctrl_wxd),
    .io_rm(fpu_io_rm),
    .io_out_x_ready(fpu_io_out_x_ready),
    .io_out_x_valid(fpu_io_out_x_valid),
    .io_out_x_bits_wb_wxd_rd(fpu_io_out_x_bits_wb_wxd_rd),
    .io_out_x_bits_wxd(fpu_io_out_x_bits_wxd),
    .io_out_x_bits_reg_idxw(fpu_io_out_x_bits_reg_idxw),
    .io_out_x_bits_warp_id(fpu_io_out_x_bits_warp_id),
    .io_out_v_ready(fpu_io_out_v_ready),
    .io_out_v_valid(fpu_io_out_v_valid),
    .io_out_v_bits_wb_wfd_rd_0(fpu_io_out_v_bits_wb_wfd_rd_0),
    .io_out_v_bits_wb_wfd_rd_1(fpu_io_out_v_bits_wb_wfd_rd_1),
    .io_out_v_bits_wb_wfd_rd_2(fpu_io_out_v_bits_wb_wfd_rd_2),
    .io_out_v_bits_wb_wfd_rd_3(fpu_io_out_v_bits_wb_wfd_rd_3),
    .io_out_v_bits_wb_wfd_rd_4(fpu_io_out_v_bits_wb_wfd_rd_4),
    .io_out_v_bits_wb_wfd_rd_5(fpu_io_out_v_bits_wb_wfd_rd_5),
    .io_out_v_bits_wb_wfd_rd_6(fpu_io_out_v_bits_wb_wfd_rd_6),
    .io_out_v_bits_wb_wfd_rd_7(fpu_io_out_v_bits_wb_wfd_rd_7),
    .io_out_v_bits_wfd_mask_0(fpu_io_out_v_bits_wfd_mask_0),
    .io_out_v_bits_wfd_mask_1(fpu_io_out_v_bits_wfd_mask_1),
    .io_out_v_bits_wfd_mask_2(fpu_io_out_v_bits_wfd_mask_2),
    .io_out_v_bits_wfd_mask_3(fpu_io_out_v_bits_wfd_mask_3),
    .io_out_v_bits_wfd_mask_4(fpu_io_out_v_bits_wfd_mask_4),
    .io_out_v_bits_wfd_mask_5(fpu_io_out_v_bits_wfd_mask_5),
    .io_out_v_bits_wfd_mask_6(fpu_io_out_v_bits_wfd_mask_6),
    .io_out_v_bits_wfd_mask_7(fpu_io_out_v_bits_wfd_mask_7),
    .io_out_v_bits_wfd(fpu_io_out_v_bits_wfd),
    .io_out_v_bits_reg_idxw(fpu_io_out_v_bits_reg_idxw),
    .io_out_v_bits_warp_id(fpu_io_out_v_bits_warp_id)
  );
  LSUexe lsu ( // @[pipe.scala 47:17]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_lsu_req_ready(lsu_io_lsu_req_ready),
    .io_lsu_req_valid(lsu_io_lsu_req_valid),
    .io_lsu_req_bits_in1_0(lsu_io_lsu_req_bits_in1_0),
    .io_lsu_req_bits_in1_1(lsu_io_lsu_req_bits_in1_1),
    .io_lsu_req_bits_in1_2(lsu_io_lsu_req_bits_in1_2),
    .io_lsu_req_bits_in1_3(lsu_io_lsu_req_bits_in1_3),
    .io_lsu_req_bits_in1_4(lsu_io_lsu_req_bits_in1_4),
    .io_lsu_req_bits_in1_5(lsu_io_lsu_req_bits_in1_5),
    .io_lsu_req_bits_in1_6(lsu_io_lsu_req_bits_in1_6),
    .io_lsu_req_bits_in1_7(lsu_io_lsu_req_bits_in1_7),
    .io_lsu_req_bits_in2_0(lsu_io_lsu_req_bits_in2_0),
    .io_lsu_req_bits_in2_1(lsu_io_lsu_req_bits_in2_1),
    .io_lsu_req_bits_in2_2(lsu_io_lsu_req_bits_in2_2),
    .io_lsu_req_bits_in2_3(lsu_io_lsu_req_bits_in2_3),
    .io_lsu_req_bits_in2_4(lsu_io_lsu_req_bits_in2_4),
    .io_lsu_req_bits_in2_5(lsu_io_lsu_req_bits_in2_5),
    .io_lsu_req_bits_in2_6(lsu_io_lsu_req_bits_in2_6),
    .io_lsu_req_bits_in2_7(lsu_io_lsu_req_bits_in2_7),
    .io_lsu_req_bits_in3_0(lsu_io_lsu_req_bits_in3_0),
    .io_lsu_req_bits_in3_1(lsu_io_lsu_req_bits_in3_1),
    .io_lsu_req_bits_in3_2(lsu_io_lsu_req_bits_in3_2),
    .io_lsu_req_bits_in3_3(lsu_io_lsu_req_bits_in3_3),
    .io_lsu_req_bits_in3_4(lsu_io_lsu_req_bits_in3_4),
    .io_lsu_req_bits_in3_5(lsu_io_lsu_req_bits_in3_5),
    .io_lsu_req_bits_in3_6(lsu_io_lsu_req_bits_in3_6),
    .io_lsu_req_bits_in3_7(lsu_io_lsu_req_bits_in3_7),
    .io_lsu_req_bits_mask_0(lsu_io_lsu_req_bits_mask_0),
    .io_lsu_req_bits_mask_1(lsu_io_lsu_req_bits_mask_1),
    .io_lsu_req_bits_mask_2(lsu_io_lsu_req_bits_mask_2),
    .io_lsu_req_bits_mask_3(lsu_io_lsu_req_bits_mask_3),
    .io_lsu_req_bits_mask_4(lsu_io_lsu_req_bits_mask_4),
    .io_lsu_req_bits_mask_5(lsu_io_lsu_req_bits_mask_5),
    .io_lsu_req_bits_mask_6(lsu_io_lsu_req_bits_mask_6),
    .io_lsu_req_bits_mask_7(lsu_io_lsu_req_bits_mask_7),
    .io_lsu_req_bits_ctrl_inst(lsu_io_lsu_req_bits_ctrl_inst),
    .io_lsu_req_bits_ctrl_wid(lsu_io_lsu_req_bits_ctrl_wid),
    .io_lsu_req_bits_ctrl_fp(lsu_io_lsu_req_bits_ctrl_fp),
    .io_lsu_req_bits_ctrl_branch(lsu_io_lsu_req_bits_ctrl_branch),
    .io_lsu_req_bits_ctrl_simt_stack(lsu_io_lsu_req_bits_ctrl_simt_stack),
    .io_lsu_req_bits_ctrl_simt_stack_op(lsu_io_lsu_req_bits_ctrl_simt_stack_op),
    .io_lsu_req_bits_ctrl_barrier(lsu_io_lsu_req_bits_ctrl_barrier),
    .io_lsu_req_bits_ctrl_csr(lsu_io_lsu_req_bits_ctrl_csr),
    .io_lsu_req_bits_ctrl_reverse(lsu_io_lsu_req_bits_ctrl_reverse),
    .io_lsu_req_bits_ctrl_isvec(lsu_io_lsu_req_bits_ctrl_isvec),
    .io_lsu_req_bits_ctrl_mem_unsigned(lsu_io_lsu_req_bits_ctrl_mem_unsigned),
    .io_lsu_req_bits_ctrl_alu_fn(lsu_io_lsu_req_bits_ctrl_alu_fn),
    .io_lsu_req_bits_ctrl_mem(lsu_io_lsu_req_bits_ctrl_mem),
    .io_lsu_req_bits_ctrl_mem_cmd(lsu_io_lsu_req_bits_ctrl_mem_cmd),
    .io_lsu_req_bits_ctrl_mop(lsu_io_lsu_req_bits_ctrl_mop),
    .io_lsu_req_bits_ctrl_reg_idxw(lsu_io_lsu_req_bits_ctrl_reg_idxw),
    .io_lsu_req_bits_ctrl_wfd(lsu_io_lsu_req_bits_ctrl_wfd),
    .io_lsu_req_bits_ctrl_fence(lsu_io_lsu_req_bits_ctrl_fence),
    .io_lsu_req_bits_ctrl_sfu(lsu_io_lsu_req_bits_ctrl_sfu),
    .io_lsu_req_bits_ctrl_readmask(lsu_io_lsu_req_bits_ctrl_readmask),
    .io_lsu_req_bits_ctrl_writemask(lsu_io_lsu_req_bits_ctrl_writemask),
    .io_lsu_req_bits_ctrl_wxd(lsu_io_lsu_req_bits_ctrl_wxd),
    .io_lsu_req_bits_ctrl_pc(lsu_io_lsu_req_bits_ctrl_pc),
    .io_dcache_rsp_ready(lsu_io_dcache_rsp_ready),
    .io_dcache_rsp_valid(lsu_io_dcache_rsp_valid),
    .io_dcache_rsp_bits_instrId(lsu_io_dcache_rsp_bits_instrId),
    .io_dcache_rsp_bits_data_0(lsu_io_dcache_rsp_bits_data_0),
    .io_dcache_rsp_bits_data_1(lsu_io_dcache_rsp_bits_data_1),
    .io_dcache_rsp_bits_data_2(lsu_io_dcache_rsp_bits_data_2),
    .io_dcache_rsp_bits_data_3(lsu_io_dcache_rsp_bits_data_3),
    .io_dcache_rsp_bits_data_4(lsu_io_dcache_rsp_bits_data_4),
    .io_dcache_rsp_bits_data_5(lsu_io_dcache_rsp_bits_data_5),
    .io_dcache_rsp_bits_data_6(lsu_io_dcache_rsp_bits_data_6),
    .io_dcache_rsp_bits_data_7(lsu_io_dcache_rsp_bits_data_7),
    .io_dcache_rsp_bits_activeMask_0(lsu_io_dcache_rsp_bits_activeMask_0),
    .io_dcache_rsp_bits_activeMask_1(lsu_io_dcache_rsp_bits_activeMask_1),
    .io_dcache_rsp_bits_activeMask_2(lsu_io_dcache_rsp_bits_activeMask_2),
    .io_dcache_rsp_bits_activeMask_3(lsu_io_dcache_rsp_bits_activeMask_3),
    .io_dcache_rsp_bits_activeMask_4(lsu_io_dcache_rsp_bits_activeMask_4),
    .io_dcache_rsp_bits_activeMask_5(lsu_io_dcache_rsp_bits_activeMask_5),
    .io_dcache_rsp_bits_activeMask_6(lsu_io_dcache_rsp_bits_activeMask_6),
    .io_dcache_rsp_bits_activeMask_7(lsu_io_dcache_rsp_bits_activeMask_7),
    .io_lsu_rsp_ready(lsu_io_lsu_rsp_ready),
    .io_lsu_rsp_valid(lsu_io_lsu_rsp_valid),
    .io_lsu_rsp_bits_tag_warp_id(lsu_io_lsu_rsp_bits_tag_warp_id),
    .io_lsu_rsp_bits_tag_wfd(lsu_io_lsu_rsp_bits_tag_wfd),
    .io_lsu_rsp_bits_tag_wxd(lsu_io_lsu_rsp_bits_tag_wxd),
    .io_lsu_rsp_bits_tag_reg_idxw(lsu_io_lsu_rsp_bits_tag_reg_idxw),
    .io_lsu_rsp_bits_tag_mask_0(lsu_io_lsu_rsp_bits_tag_mask_0),
    .io_lsu_rsp_bits_tag_mask_1(lsu_io_lsu_rsp_bits_tag_mask_1),
    .io_lsu_rsp_bits_tag_mask_2(lsu_io_lsu_rsp_bits_tag_mask_2),
    .io_lsu_rsp_bits_tag_mask_3(lsu_io_lsu_rsp_bits_tag_mask_3),
    .io_lsu_rsp_bits_tag_mask_4(lsu_io_lsu_rsp_bits_tag_mask_4),
    .io_lsu_rsp_bits_tag_mask_5(lsu_io_lsu_rsp_bits_tag_mask_5),
    .io_lsu_rsp_bits_tag_mask_6(lsu_io_lsu_rsp_bits_tag_mask_6),
    .io_lsu_rsp_bits_tag_mask_7(lsu_io_lsu_rsp_bits_tag_mask_7),
    .io_lsu_rsp_bits_tag_isWrite(lsu_io_lsu_rsp_bits_tag_isWrite),
    .io_lsu_rsp_bits_data_0(lsu_io_lsu_rsp_bits_data_0),
    .io_lsu_rsp_bits_data_1(lsu_io_lsu_rsp_bits_data_1),
    .io_lsu_rsp_bits_data_2(lsu_io_lsu_rsp_bits_data_2),
    .io_lsu_rsp_bits_data_3(lsu_io_lsu_rsp_bits_data_3),
    .io_lsu_rsp_bits_data_4(lsu_io_lsu_rsp_bits_data_4),
    .io_lsu_rsp_bits_data_5(lsu_io_lsu_rsp_bits_data_5),
    .io_lsu_rsp_bits_data_6(lsu_io_lsu_rsp_bits_data_6),
    .io_lsu_rsp_bits_data_7(lsu_io_lsu_rsp_bits_data_7),
    .io_dcache_req_ready(lsu_io_dcache_req_ready),
    .io_dcache_req_valid(lsu_io_dcache_req_valid),
    .io_dcache_req_bits_instrId(lsu_io_dcache_req_bits_instrId),
    .io_dcache_req_bits_isWrite(lsu_io_dcache_req_bits_isWrite),
    .io_dcache_req_bits_tag(lsu_io_dcache_req_bits_tag),
    .io_dcache_req_bits_setIdx(lsu_io_dcache_req_bits_setIdx),
    .io_dcache_req_bits_perLaneAddr_0_activeMask(lsu_io_dcache_req_bits_perLaneAddr_0_activeMask),
    .io_dcache_req_bits_perLaneAddr_0_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_0_blockOffset),
    .io_dcache_req_bits_perLaneAddr_1_activeMask(lsu_io_dcache_req_bits_perLaneAddr_1_activeMask),
    .io_dcache_req_bits_perLaneAddr_1_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_1_blockOffset),
    .io_dcache_req_bits_perLaneAddr_2_activeMask(lsu_io_dcache_req_bits_perLaneAddr_2_activeMask),
    .io_dcache_req_bits_perLaneAddr_2_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_2_blockOffset),
    .io_dcache_req_bits_perLaneAddr_3_activeMask(lsu_io_dcache_req_bits_perLaneAddr_3_activeMask),
    .io_dcache_req_bits_perLaneAddr_3_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_3_blockOffset),
    .io_dcache_req_bits_perLaneAddr_4_activeMask(lsu_io_dcache_req_bits_perLaneAddr_4_activeMask),
    .io_dcache_req_bits_perLaneAddr_4_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_4_blockOffset),
    .io_dcache_req_bits_perLaneAddr_5_activeMask(lsu_io_dcache_req_bits_perLaneAddr_5_activeMask),
    .io_dcache_req_bits_perLaneAddr_5_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_5_blockOffset),
    .io_dcache_req_bits_perLaneAddr_6_activeMask(lsu_io_dcache_req_bits_perLaneAddr_6_activeMask),
    .io_dcache_req_bits_perLaneAddr_6_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_6_blockOffset),
    .io_dcache_req_bits_perLaneAddr_7_activeMask(lsu_io_dcache_req_bits_perLaneAddr_7_activeMask),
    .io_dcache_req_bits_perLaneAddr_7_blockOffset(lsu_io_dcache_req_bits_perLaneAddr_7_blockOffset),
    .io_dcache_req_bits_data_0(lsu_io_dcache_req_bits_data_0),
    .io_dcache_req_bits_data_1(lsu_io_dcache_req_bits_data_1),
    .io_dcache_req_bits_data_2(lsu_io_dcache_req_bits_data_2),
    .io_dcache_req_bits_data_3(lsu_io_dcache_req_bits_data_3),
    .io_dcache_req_bits_data_4(lsu_io_dcache_req_bits_data_4),
    .io_dcache_req_bits_data_5(lsu_io_dcache_req_bits_data_5),
    .io_dcache_req_bits_data_6(lsu_io_dcache_req_bits_data_6),
    .io_dcache_req_bits_data_7(lsu_io_dcache_req_bits_data_7),
    .io_shared_req_ready(lsu_io_shared_req_ready),
    .io_shared_req_valid(lsu_io_shared_req_valid),
    .io_shared_req_bits_instrId(lsu_io_shared_req_bits_instrId),
    .io_shared_req_bits_isWrite(lsu_io_shared_req_bits_isWrite),
    .io_shared_req_bits_setIdx(lsu_io_shared_req_bits_setIdx),
    .io_shared_req_bits_perLaneAddr_0_activeMask(lsu_io_shared_req_bits_perLaneAddr_0_activeMask),
    .io_shared_req_bits_perLaneAddr_0_blockOffset(lsu_io_shared_req_bits_perLaneAddr_0_blockOffset),
    .io_shared_req_bits_perLaneAddr_1_activeMask(lsu_io_shared_req_bits_perLaneAddr_1_activeMask),
    .io_shared_req_bits_perLaneAddr_1_blockOffset(lsu_io_shared_req_bits_perLaneAddr_1_blockOffset),
    .io_shared_req_bits_perLaneAddr_2_activeMask(lsu_io_shared_req_bits_perLaneAddr_2_activeMask),
    .io_shared_req_bits_perLaneAddr_2_blockOffset(lsu_io_shared_req_bits_perLaneAddr_2_blockOffset),
    .io_shared_req_bits_perLaneAddr_3_activeMask(lsu_io_shared_req_bits_perLaneAddr_3_activeMask),
    .io_shared_req_bits_perLaneAddr_3_blockOffset(lsu_io_shared_req_bits_perLaneAddr_3_blockOffset),
    .io_shared_req_bits_perLaneAddr_4_activeMask(lsu_io_shared_req_bits_perLaneAddr_4_activeMask),
    .io_shared_req_bits_perLaneAddr_4_blockOffset(lsu_io_shared_req_bits_perLaneAddr_4_blockOffset),
    .io_shared_req_bits_perLaneAddr_5_activeMask(lsu_io_shared_req_bits_perLaneAddr_5_activeMask),
    .io_shared_req_bits_perLaneAddr_5_blockOffset(lsu_io_shared_req_bits_perLaneAddr_5_blockOffset),
    .io_shared_req_bits_perLaneAddr_6_activeMask(lsu_io_shared_req_bits_perLaneAddr_6_activeMask),
    .io_shared_req_bits_perLaneAddr_6_blockOffset(lsu_io_shared_req_bits_perLaneAddr_6_blockOffset),
    .io_shared_req_bits_perLaneAddr_7_activeMask(lsu_io_shared_req_bits_perLaneAddr_7_activeMask),
    .io_shared_req_bits_perLaneAddr_7_blockOffset(lsu_io_shared_req_bits_perLaneAddr_7_blockOffset),
    .io_shared_req_bits_data_0(lsu_io_shared_req_bits_data_0),
    .io_shared_req_bits_data_1(lsu_io_shared_req_bits_data_1),
    .io_shared_req_bits_data_2(lsu_io_shared_req_bits_data_2),
    .io_shared_req_bits_data_3(lsu_io_shared_req_bits_data_3),
    .io_shared_req_bits_data_4(lsu_io_shared_req_bits_data_4),
    .io_shared_req_bits_data_5(lsu_io_shared_req_bits_data_5),
    .io_shared_req_bits_data_6(lsu_io_shared_req_bits_data_6),
    .io_shared_req_bits_data_7(lsu_io_shared_req_bits_data_7),
    .io_shared_rsp_ready(lsu_io_shared_rsp_ready),
    .io_shared_rsp_valid(lsu_io_shared_rsp_valid),
    .io_shared_rsp_bits_instrId(lsu_io_shared_rsp_bits_instrId),
    .io_shared_rsp_bits_data_0(lsu_io_shared_rsp_bits_data_0),
    .io_shared_rsp_bits_data_1(lsu_io_shared_rsp_bits_data_1),
    .io_shared_rsp_bits_data_2(lsu_io_shared_rsp_bits_data_2),
    .io_shared_rsp_bits_data_3(lsu_io_shared_rsp_bits_data_3),
    .io_shared_rsp_bits_data_4(lsu_io_shared_rsp_bits_data_4),
    .io_shared_rsp_bits_data_5(lsu_io_shared_rsp_bits_data_5),
    .io_shared_rsp_bits_data_6(lsu_io_shared_rsp_bits_data_6),
    .io_shared_rsp_bits_data_7(lsu_io_shared_rsp_bits_data_7),
    .io_shared_rsp_bits_activeMask_0(lsu_io_shared_rsp_bits_activeMask_0),
    .io_shared_rsp_bits_activeMask_1(lsu_io_shared_rsp_bits_activeMask_1),
    .io_shared_rsp_bits_activeMask_2(lsu_io_shared_rsp_bits_activeMask_2),
    .io_shared_rsp_bits_activeMask_3(lsu_io_shared_rsp_bits_activeMask_3),
    .io_shared_rsp_bits_activeMask_4(lsu_io_shared_rsp_bits_activeMask_4),
    .io_shared_rsp_bits_activeMask_5(lsu_io_shared_rsp_bits_activeMask_5),
    .io_shared_rsp_bits_activeMask_6(lsu_io_shared_rsp_bits_activeMask_6),
    .io_shared_rsp_bits_activeMask_7(lsu_io_shared_rsp_bits_activeMask_7),
    .io_fence_end(lsu_io_fence_end)
  );
  SFUexe sfu ( // @[pipe.scala 48:17]
    .clock(sfu_clock),
    .reset(sfu_reset),
    .io_in_ready(sfu_io_in_ready),
    .io_in_valid(sfu_io_in_valid),
    .io_in_bits_in1_0(sfu_io_in_bits_in1_0),
    .io_in_bits_in1_1(sfu_io_in_bits_in1_1),
    .io_in_bits_in1_2(sfu_io_in_bits_in1_2),
    .io_in_bits_in1_3(sfu_io_in_bits_in1_3),
    .io_in_bits_in1_4(sfu_io_in_bits_in1_4),
    .io_in_bits_in1_5(sfu_io_in_bits_in1_5),
    .io_in_bits_in1_6(sfu_io_in_bits_in1_6),
    .io_in_bits_in1_7(sfu_io_in_bits_in1_7),
    .io_in_bits_in2_0(sfu_io_in_bits_in2_0),
    .io_in_bits_in2_1(sfu_io_in_bits_in2_1),
    .io_in_bits_in2_2(sfu_io_in_bits_in2_2),
    .io_in_bits_in2_3(sfu_io_in_bits_in2_3),
    .io_in_bits_in2_4(sfu_io_in_bits_in2_4),
    .io_in_bits_in2_5(sfu_io_in_bits_in2_5),
    .io_in_bits_in2_6(sfu_io_in_bits_in2_6),
    .io_in_bits_in2_7(sfu_io_in_bits_in2_7),
    .io_in_bits_mask_0(sfu_io_in_bits_mask_0),
    .io_in_bits_mask_1(sfu_io_in_bits_mask_1),
    .io_in_bits_mask_2(sfu_io_in_bits_mask_2),
    .io_in_bits_mask_3(sfu_io_in_bits_mask_3),
    .io_in_bits_mask_4(sfu_io_in_bits_mask_4),
    .io_in_bits_mask_5(sfu_io_in_bits_mask_5),
    .io_in_bits_mask_6(sfu_io_in_bits_mask_6),
    .io_in_bits_mask_7(sfu_io_in_bits_mask_7),
    .io_in_bits_ctrl_wid(sfu_io_in_bits_ctrl_wid),
    .io_in_bits_ctrl_fp(sfu_io_in_bits_ctrl_fp),
    .io_in_bits_ctrl_reverse(sfu_io_in_bits_ctrl_reverse),
    .io_in_bits_ctrl_isvec(sfu_io_in_bits_ctrl_isvec),
    .io_in_bits_ctrl_alu_fn(sfu_io_in_bits_ctrl_alu_fn),
    .io_in_bits_ctrl_reg_idxw(sfu_io_in_bits_ctrl_reg_idxw),
    .io_in_bits_ctrl_wfd(sfu_io_in_bits_ctrl_wfd),
    .io_in_bits_ctrl_wxd(sfu_io_in_bits_ctrl_wxd),
    .io_rm(sfu_io_rm),
    .io_out_x_ready(sfu_io_out_x_ready),
    .io_out_x_valid(sfu_io_out_x_valid),
    .io_out_x_bits_wb_wxd_rd(sfu_io_out_x_bits_wb_wxd_rd),
    .io_out_x_bits_wxd(sfu_io_out_x_bits_wxd),
    .io_out_x_bits_reg_idxw(sfu_io_out_x_bits_reg_idxw),
    .io_out_x_bits_warp_id(sfu_io_out_x_bits_warp_id),
    .io_out_v_ready(sfu_io_out_v_ready),
    .io_out_v_valid(sfu_io_out_v_valid),
    .io_out_v_bits_wb_wfd_rd_0(sfu_io_out_v_bits_wb_wfd_rd_0),
    .io_out_v_bits_wb_wfd_rd_1(sfu_io_out_v_bits_wb_wfd_rd_1),
    .io_out_v_bits_wb_wfd_rd_2(sfu_io_out_v_bits_wb_wfd_rd_2),
    .io_out_v_bits_wb_wfd_rd_3(sfu_io_out_v_bits_wb_wfd_rd_3),
    .io_out_v_bits_wb_wfd_rd_4(sfu_io_out_v_bits_wb_wfd_rd_4),
    .io_out_v_bits_wb_wfd_rd_5(sfu_io_out_v_bits_wb_wfd_rd_5),
    .io_out_v_bits_wb_wfd_rd_6(sfu_io_out_v_bits_wb_wfd_rd_6),
    .io_out_v_bits_wb_wfd_rd_7(sfu_io_out_v_bits_wb_wfd_rd_7),
    .io_out_v_bits_wfd_mask_0(sfu_io_out_v_bits_wfd_mask_0),
    .io_out_v_bits_wfd_mask_1(sfu_io_out_v_bits_wfd_mask_1),
    .io_out_v_bits_wfd_mask_2(sfu_io_out_v_bits_wfd_mask_2),
    .io_out_v_bits_wfd_mask_3(sfu_io_out_v_bits_wfd_mask_3),
    .io_out_v_bits_wfd_mask_4(sfu_io_out_v_bits_wfd_mask_4),
    .io_out_v_bits_wfd_mask_5(sfu_io_out_v_bits_wfd_mask_5),
    .io_out_v_bits_wfd_mask_6(sfu_io_out_v_bits_wfd_mask_6),
    .io_out_v_bits_wfd_mask_7(sfu_io_out_v_bits_wfd_mask_7),
    .io_out_v_bits_wfd(sfu_io_out_v_bits_wfd),
    .io_out_v_bits_reg_idxw(sfu_io_out_v_bits_reg_idxw),
    .io_out_v_bits_warp_id(sfu_io_out_v_bits_warp_id)
  );
  LSU2WB lsu2wb ( // @[pipe.scala 49:20]
    .io_lsu_rsp_ready(lsu2wb_io_lsu_rsp_ready),
    .io_lsu_rsp_valid(lsu2wb_io_lsu_rsp_valid),
    .io_lsu_rsp_bits_tag_warp_id(lsu2wb_io_lsu_rsp_bits_tag_warp_id),
    .io_lsu_rsp_bits_tag_wfd(lsu2wb_io_lsu_rsp_bits_tag_wfd),
    .io_lsu_rsp_bits_tag_wxd(lsu2wb_io_lsu_rsp_bits_tag_wxd),
    .io_lsu_rsp_bits_tag_reg_idxw(lsu2wb_io_lsu_rsp_bits_tag_reg_idxw),
    .io_lsu_rsp_bits_tag_mask_0(lsu2wb_io_lsu_rsp_bits_tag_mask_0),
    .io_lsu_rsp_bits_tag_mask_1(lsu2wb_io_lsu_rsp_bits_tag_mask_1),
    .io_lsu_rsp_bits_tag_mask_2(lsu2wb_io_lsu_rsp_bits_tag_mask_2),
    .io_lsu_rsp_bits_tag_mask_3(lsu2wb_io_lsu_rsp_bits_tag_mask_3),
    .io_lsu_rsp_bits_tag_mask_4(lsu2wb_io_lsu_rsp_bits_tag_mask_4),
    .io_lsu_rsp_bits_tag_mask_5(lsu2wb_io_lsu_rsp_bits_tag_mask_5),
    .io_lsu_rsp_bits_tag_mask_6(lsu2wb_io_lsu_rsp_bits_tag_mask_6),
    .io_lsu_rsp_bits_tag_mask_7(lsu2wb_io_lsu_rsp_bits_tag_mask_7),
    .io_lsu_rsp_bits_tag_isWrite(lsu2wb_io_lsu_rsp_bits_tag_isWrite),
    .io_lsu_rsp_bits_data_0(lsu2wb_io_lsu_rsp_bits_data_0),
    .io_lsu_rsp_bits_data_1(lsu2wb_io_lsu_rsp_bits_data_1),
    .io_lsu_rsp_bits_data_2(lsu2wb_io_lsu_rsp_bits_data_2),
    .io_lsu_rsp_bits_data_3(lsu2wb_io_lsu_rsp_bits_data_3),
    .io_lsu_rsp_bits_data_4(lsu2wb_io_lsu_rsp_bits_data_4),
    .io_lsu_rsp_bits_data_5(lsu2wb_io_lsu_rsp_bits_data_5),
    .io_lsu_rsp_bits_data_6(lsu2wb_io_lsu_rsp_bits_data_6),
    .io_lsu_rsp_bits_data_7(lsu2wb_io_lsu_rsp_bits_data_7),
    .io_out_x_ready(lsu2wb_io_out_x_ready),
    .io_out_x_valid(lsu2wb_io_out_x_valid),
    .io_out_x_bits_wb_wxd_rd(lsu2wb_io_out_x_bits_wb_wxd_rd),
    .io_out_x_bits_wxd(lsu2wb_io_out_x_bits_wxd),
    .io_out_x_bits_reg_idxw(lsu2wb_io_out_x_bits_reg_idxw),
    .io_out_x_bits_warp_id(lsu2wb_io_out_x_bits_warp_id),
    .io_out_v_ready(lsu2wb_io_out_v_ready),
    .io_out_v_valid(lsu2wb_io_out_v_valid),
    .io_out_v_bits_wb_wfd_rd_0(lsu2wb_io_out_v_bits_wb_wfd_rd_0),
    .io_out_v_bits_wb_wfd_rd_1(lsu2wb_io_out_v_bits_wb_wfd_rd_1),
    .io_out_v_bits_wb_wfd_rd_2(lsu2wb_io_out_v_bits_wb_wfd_rd_2),
    .io_out_v_bits_wb_wfd_rd_3(lsu2wb_io_out_v_bits_wb_wfd_rd_3),
    .io_out_v_bits_wb_wfd_rd_4(lsu2wb_io_out_v_bits_wb_wfd_rd_4),
    .io_out_v_bits_wb_wfd_rd_5(lsu2wb_io_out_v_bits_wb_wfd_rd_5),
    .io_out_v_bits_wb_wfd_rd_6(lsu2wb_io_out_v_bits_wb_wfd_rd_6),
    .io_out_v_bits_wb_wfd_rd_7(lsu2wb_io_out_v_bits_wb_wfd_rd_7),
    .io_out_v_bits_wfd_mask_0(lsu2wb_io_out_v_bits_wfd_mask_0),
    .io_out_v_bits_wfd_mask_1(lsu2wb_io_out_v_bits_wfd_mask_1),
    .io_out_v_bits_wfd_mask_2(lsu2wb_io_out_v_bits_wfd_mask_2),
    .io_out_v_bits_wfd_mask_3(lsu2wb_io_out_v_bits_wfd_mask_3),
    .io_out_v_bits_wfd_mask_4(lsu2wb_io_out_v_bits_wfd_mask_4),
    .io_out_v_bits_wfd_mask_5(lsu2wb_io_out_v_bits_wfd_mask_5),
    .io_out_v_bits_wfd_mask_6(lsu2wb_io_out_v_bits_wfd_mask_6),
    .io_out_v_bits_wfd_mask_7(lsu2wb_io_out_v_bits_wfd_mask_7),
    .io_out_v_bits_wfd(lsu2wb_io_out_v_bits_wfd),
    .io_out_v_bits_reg_idxw(lsu2wb_io_out_v_bits_reg_idxw),
    .io_out_v_bits_warp_id(lsu2wb_io_out_v_bits_warp_id)
  );
  Writeback wb ( // @[pipe.scala 50:16]
    .io_out_v_ready(wb_io_out_v_ready),
    .io_out_v_valid(wb_io_out_v_valid),
    .io_out_v_bits_wb_wfd_rd_0(wb_io_out_v_bits_wb_wfd_rd_0),
    .io_out_v_bits_wb_wfd_rd_1(wb_io_out_v_bits_wb_wfd_rd_1),
    .io_out_v_bits_wb_wfd_rd_2(wb_io_out_v_bits_wb_wfd_rd_2),
    .io_out_v_bits_wb_wfd_rd_3(wb_io_out_v_bits_wb_wfd_rd_3),
    .io_out_v_bits_wb_wfd_rd_4(wb_io_out_v_bits_wb_wfd_rd_4),
    .io_out_v_bits_wb_wfd_rd_5(wb_io_out_v_bits_wb_wfd_rd_5),
    .io_out_v_bits_wb_wfd_rd_6(wb_io_out_v_bits_wb_wfd_rd_6),
    .io_out_v_bits_wb_wfd_rd_7(wb_io_out_v_bits_wb_wfd_rd_7),
    .io_out_v_bits_wfd_mask_0(wb_io_out_v_bits_wfd_mask_0),
    .io_out_v_bits_wfd_mask_1(wb_io_out_v_bits_wfd_mask_1),
    .io_out_v_bits_wfd_mask_2(wb_io_out_v_bits_wfd_mask_2),
    .io_out_v_bits_wfd_mask_3(wb_io_out_v_bits_wfd_mask_3),
    .io_out_v_bits_wfd_mask_4(wb_io_out_v_bits_wfd_mask_4),
    .io_out_v_bits_wfd_mask_5(wb_io_out_v_bits_wfd_mask_5),
    .io_out_v_bits_wfd_mask_6(wb_io_out_v_bits_wfd_mask_6),
    .io_out_v_bits_wfd_mask_7(wb_io_out_v_bits_wfd_mask_7),
    .io_out_v_bits_wfd(wb_io_out_v_bits_wfd),
    .io_out_v_bits_reg_idxw(wb_io_out_v_bits_reg_idxw),
    .io_out_v_bits_warp_id(wb_io_out_v_bits_warp_id),
    .io_out_x_ready(wb_io_out_x_ready),
    .io_out_x_valid(wb_io_out_x_valid),
    .io_out_x_bits_wb_wxd_rd(wb_io_out_x_bits_wb_wxd_rd),
    .io_out_x_bits_wxd(wb_io_out_x_bits_wxd),
    .io_out_x_bits_reg_idxw(wb_io_out_x_bits_reg_idxw),
    .io_out_x_bits_warp_id(wb_io_out_x_bits_warp_id),
    .io_in_x_0_valid(wb_io_in_x_0_valid),
    .io_in_x_0_bits_wb_wxd_rd(wb_io_in_x_0_bits_wb_wxd_rd),
    .io_in_x_0_bits_wxd(wb_io_in_x_0_bits_wxd),
    .io_in_x_0_bits_reg_idxw(wb_io_in_x_0_bits_reg_idxw),
    .io_in_x_0_bits_warp_id(wb_io_in_x_0_bits_warp_id),
    .io_in_x_1_ready(wb_io_in_x_1_ready),
    .io_in_x_1_valid(wb_io_in_x_1_valid),
    .io_in_x_1_bits_wb_wxd_rd(wb_io_in_x_1_bits_wb_wxd_rd),
    .io_in_x_1_bits_wxd(wb_io_in_x_1_bits_wxd),
    .io_in_x_1_bits_reg_idxw(wb_io_in_x_1_bits_reg_idxw),
    .io_in_x_1_bits_warp_id(wb_io_in_x_1_bits_warp_id),
    .io_in_x_2_ready(wb_io_in_x_2_ready),
    .io_in_x_2_valid(wb_io_in_x_2_valid),
    .io_in_x_2_bits_wb_wxd_rd(wb_io_in_x_2_bits_wb_wxd_rd),
    .io_in_x_2_bits_wxd(wb_io_in_x_2_bits_wxd),
    .io_in_x_2_bits_reg_idxw(wb_io_in_x_2_bits_reg_idxw),
    .io_in_x_2_bits_warp_id(wb_io_in_x_2_bits_warp_id),
    .io_in_x_3_ready(wb_io_in_x_3_ready),
    .io_in_x_3_valid(wb_io_in_x_3_valid),
    .io_in_x_3_bits_wb_wxd_rd(wb_io_in_x_3_bits_wb_wxd_rd),
    .io_in_x_3_bits_wxd(wb_io_in_x_3_bits_wxd),
    .io_in_x_3_bits_reg_idxw(wb_io_in_x_3_bits_reg_idxw),
    .io_in_x_3_bits_warp_id(wb_io_in_x_3_bits_warp_id),
    .io_in_x_4_ready(wb_io_in_x_4_ready),
    .io_in_x_4_valid(wb_io_in_x_4_valid),
    .io_in_x_4_bits_wb_wxd_rd(wb_io_in_x_4_bits_wb_wxd_rd),
    .io_in_x_4_bits_wxd(wb_io_in_x_4_bits_wxd),
    .io_in_x_4_bits_reg_idxw(wb_io_in_x_4_bits_reg_idxw),
    .io_in_x_4_bits_warp_id(wb_io_in_x_4_bits_warp_id),
    .io_in_v_0_valid(wb_io_in_v_0_valid),
    .io_in_v_0_bits_wb_wfd_rd_0(wb_io_in_v_0_bits_wb_wfd_rd_0),
    .io_in_v_0_bits_wb_wfd_rd_1(wb_io_in_v_0_bits_wb_wfd_rd_1),
    .io_in_v_0_bits_wb_wfd_rd_2(wb_io_in_v_0_bits_wb_wfd_rd_2),
    .io_in_v_0_bits_wb_wfd_rd_3(wb_io_in_v_0_bits_wb_wfd_rd_3),
    .io_in_v_0_bits_wb_wfd_rd_4(wb_io_in_v_0_bits_wb_wfd_rd_4),
    .io_in_v_0_bits_wb_wfd_rd_5(wb_io_in_v_0_bits_wb_wfd_rd_5),
    .io_in_v_0_bits_wb_wfd_rd_6(wb_io_in_v_0_bits_wb_wfd_rd_6),
    .io_in_v_0_bits_wb_wfd_rd_7(wb_io_in_v_0_bits_wb_wfd_rd_7),
    .io_in_v_0_bits_wfd_mask_0(wb_io_in_v_0_bits_wfd_mask_0),
    .io_in_v_0_bits_wfd_mask_1(wb_io_in_v_0_bits_wfd_mask_1),
    .io_in_v_0_bits_wfd_mask_2(wb_io_in_v_0_bits_wfd_mask_2),
    .io_in_v_0_bits_wfd_mask_3(wb_io_in_v_0_bits_wfd_mask_3),
    .io_in_v_0_bits_wfd_mask_4(wb_io_in_v_0_bits_wfd_mask_4),
    .io_in_v_0_bits_wfd_mask_5(wb_io_in_v_0_bits_wfd_mask_5),
    .io_in_v_0_bits_wfd_mask_6(wb_io_in_v_0_bits_wfd_mask_6),
    .io_in_v_0_bits_wfd_mask_7(wb_io_in_v_0_bits_wfd_mask_7),
    .io_in_v_0_bits_wfd(wb_io_in_v_0_bits_wfd),
    .io_in_v_0_bits_reg_idxw(wb_io_in_v_0_bits_reg_idxw),
    .io_in_v_0_bits_warp_id(wb_io_in_v_0_bits_warp_id),
    .io_in_v_1_ready(wb_io_in_v_1_ready),
    .io_in_v_1_valid(wb_io_in_v_1_valid),
    .io_in_v_1_bits_wb_wfd_rd_0(wb_io_in_v_1_bits_wb_wfd_rd_0),
    .io_in_v_1_bits_wb_wfd_rd_1(wb_io_in_v_1_bits_wb_wfd_rd_1),
    .io_in_v_1_bits_wb_wfd_rd_2(wb_io_in_v_1_bits_wb_wfd_rd_2),
    .io_in_v_1_bits_wb_wfd_rd_3(wb_io_in_v_1_bits_wb_wfd_rd_3),
    .io_in_v_1_bits_wb_wfd_rd_4(wb_io_in_v_1_bits_wb_wfd_rd_4),
    .io_in_v_1_bits_wb_wfd_rd_5(wb_io_in_v_1_bits_wb_wfd_rd_5),
    .io_in_v_1_bits_wb_wfd_rd_6(wb_io_in_v_1_bits_wb_wfd_rd_6),
    .io_in_v_1_bits_wb_wfd_rd_7(wb_io_in_v_1_bits_wb_wfd_rd_7),
    .io_in_v_1_bits_wfd_mask_0(wb_io_in_v_1_bits_wfd_mask_0),
    .io_in_v_1_bits_wfd_mask_1(wb_io_in_v_1_bits_wfd_mask_1),
    .io_in_v_1_bits_wfd_mask_2(wb_io_in_v_1_bits_wfd_mask_2),
    .io_in_v_1_bits_wfd_mask_3(wb_io_in_v_1_bits_wfd_mask_3),
    .io_in_v_1_bits_wfd_mask_4(wb_io_in_v_1_bits_wfd_mask_4),
    .io_in_v_1_bits_wfd_mask_5(wb_io_in_v_1_bits_wfd_mask_5),
    .io_in_v_1_bits_wfd_mask_6(wb_io_in_v_1_bits_wfd_mask_6),
    .io_in_v_1_bits_wfd_mask_7(wb_io_in_v_1_bits_wfd_mask_7),
    .io_in_v_1_bits_wfd(wb_io_in_v_1_bits_wfd),
    .io_in_v_1_bits_reg_idxw(wb_io_in_v_1_bits_reg_idxw),
    .io_in_v_1_bits_warp_id(wb_io_in_v_1_bits_warp_id),
    .io_in_v_2_ready(wb_io_in_v_2_ready),
    .io_in_v_2_valid(wb_io_in_v_2_valid),
    .io_in_v_2_bits_wb_wfd_rd_0(wb_io_in_v_2_bits_wb_wfd_rd_0),
    .io_in_v_2_bits_wb_wfd_rd_1(wb_io_in_v_2_bits_wb_wfd_rd_1),
    .io_in_v_2_bits_wb_wfd_rd_2(wb_io_in_v_2_bits_wb_wfd_rd_2),
    .io_in_v_2_bits_wb_wfd_rd_3(wb_io_in_v_2_bits_wb_wfd_rd_3),
    .io_in_v_2_bits_wb_wfd_rd_4(wb_io_in_v_2_bits_wb_wfd_rd_4),
    .io_in_v_2_bits_wb_wfd_rd_5(wb_io_in_v_2_bits_wb_wfd_rd_5),
    .io_in_v_2_bits_wb_wfd_rd_6(wb_io_in_v_2_bits_wb_wfd_rd_6),
    .io_in_v_2_bits_wb_wfd_rd_7(wb_io_in_v_2_bits_wb_wfd_rd_7),
    .io_in_v_2_bits_wfd_mask_0(wb_io_in_v_2_bits_wfd_mask_0),
    .io_in_v_2_bits_wfd_mask_1(wb_io_in_v_2_bits_wfd_mask_1),
    .io_in_v_2_bits_wfd_mask_2(wb_io_in_v_2_bits_wfd_mask_2),
    .io_in_v_2_bits_wfd_mask_3(wb_io_in_v_2_bits_wfd_mask_3),
    .io_in_v_2_bits_wfd_mask_4(wb_io_in_v_2_bits_wfd_mask_4),
    .io_in_v_2_bits_wfd_mask_5(wb_io_in_v_2_bits_wfd_mask_5),
    .io_in_v_2_bits_wfd_mask_6(wb_io_in_v_2_bits_wfd_mask_6),
    .io_in_v_2_bits_wfd_mask_7(wb_io_in_v_2_bits_wfd_mask_7),
    .io_in_v_2_bits_wfd(wb_io_in_v_2_bits_wfd),
    .io_in_v_2_bits_reg_idxw(wb_io_in_v_2_bits_reg_idxw),
    .io_in_v_2_bits_warp_id(wb_io_in_v_2_bits_warp_id),
    .io_in_v_3_ready(wb_io_in_v_3_ready),
    .io_in_v_3_valid(wb_io_in_v_3_valid),
    .io_in_v_3_bits_wb_wfd_rd_0(wb_io_in_v_3_bits_wb_wfd_rd_0),
    .io_in_v_3_bits_wb_wfd_rd_1(wb_io_in_v_3_bits_wb_wfd_rd_1),
    .io_in_v_3_bits_wb_wfd_rd_2(wb_io_in_v_3_bits_wb_wfd_rd_2),
    .io_in_v_3_bits_wb_wfd_rd_3(wb_io_in_v_3_bits_wb_wfd_rd_3),
    .io_in_v_3_bits_wb_wfd_rd_4(wb_io_in_v_3_bits_wb_wfd_rd_4),
    .io_in_v_3_bits_wb_wfd_rd_5(wb_io_in_v_3_bits_wb_wfd_rd_5),
    .io_in_v_3_bits_wb_wfd_rd_6(wb_io_in_v_3_bits_wb_wfd_rd_6),
    .io_in_v_3_bits_wb_wfd_rd_7(wb_io_in_v_3_bits_wb_wfd_rd_7),
    .io_in_v_3_bits_wfd_mask_0(wb_io_in_v_3_bits_wfd_mask_0),
    .io_in_v_3_bits_wfd_mask_1(wb_io_in_v_3_bits_wfd_mask_1),
    .io_in_v_3_bits_wfd_mask_2(wb_io_in_v_3_bits_wfd_mask_2),
    .io_in_v_3_bits_wfd_mask_3(wb_io_in_v_3_bits_wfd_mask_3),
    .io_in_v_3_bits_wfd_mask_4(wb_io_in_v_3_bits_wfd_mask_4),
    .io_in_v_3_bits_wfd_mask_5(wb_io_in_v_3_bits_wfd_mask_5),
    .io_in_v_3_bits_wfd_mask_6(wb_io_in_v_3_bits_wfd_mask_6),
    .io_in_v_3_bits_wfd_mask_7(wb_io_in_v_3_bits_wfd_mask_7),
    .io_in_v_3_bits_wfd(wb_io_in_v_3_bits_wfd),
    .io_in_v_3_bits_reg_idxw(wb_io_in_v_3_bits_reg_idxw),
    .io_in_v_3_bits_warp_id(wb_io_in_v_3_bits_warp_id)
  );
  Scoreboard Scoreboard ( // @[pipe.scala 52:47]
    .clock(Scoreboard_clock),
    .reset(Scoreboard_reset),
    .io_ibuffer_if_ctrl_sel_alu2(Scoreboard_io_ibuffer_if_ctrl_sel_alu2),
    .io_ibuffer_if_ctrl_sel_alu1(Scoreboard_io_ibuffer_if_ctrl_sel_alu1),
    .io_ibuffer_if_ctrl_isvec(Scoreboard_io_ibuffer_if_ctrl_isvec),
    .io_ibuffer_if_ctrl_sel_alu3(Scoreboard_io_ibuffer_if_ctrl_sel_alu3),
    .io_ibuffer_if_ctrl_mask(Scoreboard_io_ibuffer_if_ctrl_mask),
    .io_ibuffer_if_ctrl_mem(Scoreboard_io_ibuffer_if_ctrl_mem),
    .io_ibuffer_if_ctrl_reg_idx1(Scoreboard_io_ibuffer_if_ctrl_reg_idx1),
    .io_ibuffer_if_ctrl_reg_idx2(Scoreboard_io_ibuffer_if_ctrl_reg_idx2),
    .io_ibuffer_if_ctrl_reg_idx3(Scoreboard_io_ibuffer_if_ctrl_reg_idx3),
    .io_if_ctrl_branch(Scoreboard_io_if_ctrl_branch),
    .io_if_ctrl_barrier(Scoreboard_io_if_ctrl_barrier),
    .io_if_ctrl_reg_idxw(Scoreboard_io_if_ctrl_reg_idxw),
    .io_if_ctrl_wfd(Scoreboard_io_if_ctrl_wfd),
    .io_if_ctrl_fence(Scoreboard_io_if_ctrl_fence),
    .io_if_ctrl_wxd(Scoreboard_io_if_ctrl_wxd),
    .io_wb_v_ctrl_wfd(Scoreboard_io_wb_v_ctrl_wfd),
    .io_wb_v_ctrl_reg_idxw(Scoreboard_io_wb_v_ctrl_reg_idxw),
    .io_wb_x_ctrl_wxd(Scoreboard_io_wb_x_ctrl_wxd),
    .io_wb_x_ctrl_reg_idxw(Scoreboard_io_wb_x_ctrl_reg_idxw),
    .io_if_fire(Scoreboard_io_if_fire),
    .io_br_ctrl(Scoreboard_io_br_ctrl),
    .io_fence_end(Scoreboard_io_fence_end),
    .io_wb_v_fire(Scoreboard_io_wb_v_fire),
    .io_wb_x_fire(Scoreboard_io_wb_x_fire),
    .io_delay(Scoreboard_io_delay)
  );
  Scoreboard Scoreboard_1 ( // @[pipe.scala 52:47]
    .clock(Scoreboard_1_clock),
    .reset(Scoreboard_1_reset),
    .io_ibuffer_if_ctrl_sel_alu2(Scoreboard_1_io_ibuffer_if_ctrl_sel_alu2),
    .io_ibuffer_if_ctrl_sel_alu1(Scoreboard_1_io_ibuffer_if_ctrl_sel_alu1),
    .io_ibuffer_if_ctrl_isvec(Scoreboard_1_io_ibuffer_if_ctrl_isvec),
    .io_ibuffer_if_ctrl_sel_alu3(Scoreboard_1_io_ibuffer_if_ctrl_sel_alu3),
    .io_ibuffer_if_ctrl_mask(Scoreboard_1_io_ibuffer_if_ctrl_mask),
    .io_ibuffer_if_ctrl_mem(Scoreboard_1_io_ibuffer_if_ctrl_mem),
    .io_ibuffer_if_ctrl_reg_idx1(Scoreboard_1_io_ibuffer_if_ctrl_reg_idx1),
    .io_ibuffer_if_ctrl_reg_idx2(Scoreboard_1_io_ibuffer_if_ctrl_reg_idx2),
    .io_ibuffer_if_ctrl_reg_idx3(Scoreboard_1_io_ibuffer_if_ctrl_reg_idx3),
    .io_if_ctrl_branch(Scoreboard_1_io_if_ctrl_branch),
    .io_if_ctrl_barrier(Scoreboard_1_io_if_ctrl_barrier),
    .io_if_ctrl_reg_idxw(Scoreboard_1_io_if_ctrl_reg_idxw),
    .io_if_ctrl_wfd(Scoreboard_1_io_if_ctrl_wfd),
    .io_if_ctrl_fence(Scoreboard_1_io_if_ctrl_fence),
    .io_if_ctrl_wxd(Scoreboard_1_io_if_ctrl_wxd),
    .io_wb_v_ctrl_wfd(Scoreboard_1_io_wb_v_ctrl_wfd),
    .io_wb_v_ctrl_reg_idxw(Scoreboard_1_io_wb_v_ctrl_reg_idxw),
    .io_wb_x_ctrl_wxd(Scoreboard_1_io_wb_x_ctrl_wxd),
    .io_wb_x_ctrl_reg_idxw(Scoreboard_1_io_wb_x_ctrl_reg_idxw),
    .io_if_fire(Scoreboard_1_io_if_fire),
    .io_br_ctrl(Scoreboard_1_io_br_ctrl),
    .io_fence_end(Scoreboard_1_io_fence_end),
    .io_wb_v_fire(Scoreboard_1_io_wb_v_fire),
    .io_wb_x_fire(Scoreboard_1_io_wb_x_fire),
    .io_delay(Scoreboard_1_io_delay)
  );
  Scoreboard Scoreboard_2 ( // @[pipe.scala 52:47]
    .clock(Scoreboard_2_clock),
    .reset(Scoreboard_2_reset),
    .io_ibuffer_if_ctrl_sel_alu2(Scoreboard_2_io_ibuffer_if_ctrl_sel_alu2),
    .io_ibuffer_if_ctrl_sel_alu1(Scoreboard_2_io_ibuffer_if_ctrl_sel_alu1),
    .io_ibuffer_if_ctrl_isvec(Scoreboard_2_io_ibuffer_if_ctrl_isvec),
    .io_ibuffer_if_ctrl_sel_alu3(Scoreboard_2_io_ibuffer_if_ctrl_sel_alu3),
    .io_ibuffer_if_ctrl_mask(Scoreboard_2_io_ibuffer_if_ctrl_mask),
    .io_ibuffer_if_ctrl_mem(Scoreboard_2_io_ibuffer_if_ctrl_mem),
    .io_ibuffer_if_ctrl_reg_idx1(Scoreboard_2_io_ibuffer_if_ctrl_reg_idx1),
    .io_ibuffer_if_ctrl_reg_idx2(Scoreboard_2_io_ibuffer_if_ctrl_reg_idx2),
    .io_ibuffer_if_ctrl_reg_idx3(Scoreboard_2_io_ibuffer_if_ctrl_reg_idx3),
    .io_if_ctrl_branch(Scoreboard_2_io_if_ctrl_branch),
    .io_if_ctrl_barrier(Scoreboard_2_io_if_ctrl_barrier),
    .io_if_ctrl_reg_idxw(Scoreboard_2_io_if_ctrl_reg_idxw),
    .io_if_ctrl_wfd(Scoreboard_2_io_if_ctrl_wfd),
    .io_if_ctrl_fence(Scoreboard_2_io_if_ctrl_fence),
    .io_if_ctrl_wxd(Scoreboard_2_io_if_ctrl_wxd),
    .io_wb_v_ctrl_wfd(Scoreboard_2_io_wb_v_ctrl_wfd),
    .io_wb_v_ctrl_reg_idxw(Scoreboard_2_io_wb_v_ctrl_reg_idxw),
    .io_wb_x_ctrl_wxd(Scoreboard_2_io_wb_x_ctrl_wxd),
    .io_wb_x_ctrl_reg_idxw(Scoreboard_2_io_wb_x_ctrl_reg_idxw),
    .io_if_fire(Scoreboard_2_io_if_fire),
    .io_br_ctrl(Scoreboard_2_io_br_ctrl),
    .io_fence_end(Scoreboard_2_io_fence_end),
    .io_wb_v_fire(Scoreboard_2_io_wb_v_fire),
    .io_wb_x_fire(Scoreboard_2_io_wb_x_fire),
    .io_delay(Scoreboard_2_io_delay)
  );
  Scoreboard Scoreboard_3 ( // @[pipe.scala 52:47]
    .clock(Scoreboard_3_clock),
    .reset(Scoreboard_3_reset),
    .io_ibuffer_if_ctrl_sel_alu2(Scoreboard_3_io_ibuffer_if_ctrl_sel_alu2),
    .io_ibuffer_if_ctrl_sel_alu1(Scoreboard_3_io_ibuffer_if_ctrl_sel_alu1),
    .io_ibuffer_if_ctrl_isvec(Scoreboard_3_io_ibuffer_if_ctrl_isvec),
    .io_ibuffer_if_ctrl_sel_alu3(Scoreboard_3_io_ibuffer_if_ctrl_sel_alu3),
    .io_ibuffer_if_ctrl_mask(Scoreboard_3_io_ibuffer_if_ctrl_mask),
    .io_ibuffer_if_ctrl_mem(Scoreboard_3_io_ibuffer_if_ctrl_mem),
    .io_ibuffer_if_ctrl_reg_idx1(Scoreboard_3_io_ibuffer_if_ctrl_reg_idx1),
    .io_ibuffer_if_ctrl_reg_idx2(Scoreboard_3_io_ibuffer_if_ctrl_reg_idx2),
    .io_ibuffer_if_ctrl_reg_idx3(Scoreboard_3_io_ibuffer_if_ctrl_reg_idx3),
    .io_if_ctrl_branch(Scoreboard_3_io_if_ctrl_branch),
    .io_if_ctrl_barrier(Scoreboard_3_io_if_ctrl_barrier),
    .io_if_ctrl_reg_idxw(Scoreboard_3_io_if_ctrl_reg_idxw),
    .io_if_ctrl_wfd(Scoreboard_3_io_if_ctrl_wfd),
    .io_if_ctrl_fence(Scoreboard_3_io_if_ctrl_fence),
    .io_if_ctrl_wxd(Scoreboard_3_io_if_ctrl_wxd),
    .io_wb_v_ctrl_wfd(Scoreboard_3_io_wb_v_ctrl_wfd),
    .io_wb_v_ctrl_reg_idxw(Scoreboard_3_io_wb_v_ctrl_reg_idxw),
    .io_wb_x_ctrl_wxd(Scoreboard_3_io_wb_x_ctrl_wxd),
    .io_wb_x_ctrl_reg_idxw(Scoreboard_3_io_wb_x_ctrl_reg_idxw),
    .io_if_fire(Scoreboard_3_io_if_fire),
    .io_br_ctrl(Scoreboard_3_io_br_ctrl),
    .io_fence_end(Scoreboard_3_io_fence_end),
    .io_wb_v_fire(Scoreboard_3_io_wb_v_fire),
    .io_wb_x_fire(Scoreboard_3_io_wb_x_fire),
    .io_delay(Scoreboard_3_io_delay)
  );
  instbuffer ibuffer ( // @[pipe.scala 53:21]
    .clock(ibuffer_clock),
    .reset(ibuffer_reset),
    .io_in_ready(ibuffer_io_in_ready),
    .io_in_valid(ibuffer_io_in_valid),
    .io_in_bits_inst(ibuffer_io_in_bits_inst),
    .io_in_bits_wid(ibuffer_io_in_bits_wid),
    .io_in_bits_fp(ibuffer_io_in_bits_fp),
    .io_in_bits_branch(ibuffer_io_in_bits_branch),
    .io_in_bits_simt_stack(ibuffer_io_in_bits_simt_stack),
    .io_in_bits_simt_stack_op(ibuffer_io_in_bits_simt_stack_op),
    .io_in_bits_barrier(ibuffer_io_in_bits_barrier),
    .io_in_bits_csr(ibuffer_io_in_bits_csr),
    .io_in_bits_reverse(ibuffer_io_in_bits_reverse),
    .io_in_bits_sel_alu2(ibuffer_io_in_bits_sel_alu2),
    .io_in_bits_sel_alu1(ibuffer_io_in_bits_sel_alu1),
    .io_in_bits_isvec(ibuffer_io_in_bits_isvec),
    .io_in_bits_sel_alu3(ibuffer_io_in_bits_sel_alu3),
    .io_in_bits_mask(ibuffer_io_in_bits_mask),
    .io_in_bits_sel_imm(ibuffer_io_in_bits_sel_imm),
    .io_in_bits_mem_unsigned(ibuffer_io_in_bits_mem_unsigned),
    .io_in_bits_alu_fn(ibuffer_io_in_bits_alu_fn),
    .io_in_bits_mem(ibuffer_io_in_bits_mem),
    .io_in_bits_mem_cmd(ibuffer_io_in_bits_mem_cmd),
    .io_in_bits_mop(ibuffer_io_in_bits_mop),
    .io_in_bits_reg_idx1(ibuffer_io_in_bits_reg_idx1),
    .io_in_bits_reg_idx2(ibuffer_io_in_bits_reg_idx2),
    .io_in_bits_reg_idx3(ibuffer_io_in_bits_reg_idx3),
    .io_in_bits_reg_idxw(ibuffer_io_in_bits_reg_idxw),
    .io_in_bits_wfd(ibuffer_io_in_bits_wfd),
    .io_in_bits_fence(ibuffer_io_in_bits_fence),
    .io_in_bits_sfu(ibuffer_io_in_bits_sfu),
    .io_in_bits_readmask(ibuffer_io_in_bits_readmask),
    .io_in_bits_writemask(ibuffer_io_in_bits_writemask),
    .io_in_bits_wxd(ibuffer_io_in_bits_wxd),
    .io_in_bits_pc(ibuffer_io_in_bits_pc),
    .io_flush_valid(ibuffer_io_flush_valid),
    .io_flush_bits(ibuffer_io_flush_bits),
    .io_out_0_ready(ibuffer_io_out_0_ready),
    .io_out_0_valid(ibuffer_io_out_0_valid),
    .io_out_0_bits_inst(ibuffer_io_out_0_bits_inst),
    .io_out_0_bits_wid(ibuffer_io_out_0_bits_wid),
    .io_out_0_bits_fp(ibuffer_io_out_0_bits_fp),
    .io_out_0_bits_branch(ibuffer_io_out_0_bits_branch),
    .io_out_0_bits_simt_stack(ibuffer_io_out_0_bits_simt_stack),
    .io_out_0_bits_simt_stack_op(ibuffer_io_out_0_bits_simt_stack_op),
    .io_out_0_bits_barrier(ibuffer_io_out_0_bits_barrier),
    .io_out_0_bits_csr(ibuffer_io_out_0_bits_csr),
    .io_out_0_bits_reverse(ibuffer_io_out_0_bits_reverse),
    .io_out_0_bits_sel_alu2(ibuffer_io_out_0_bits_sel_alu2),
    .io_out_0_bits_sel_alu1(ibuffer_io_out_0_bits_sel_alu1),
    .io_out_0_bits_isvec(ibuffer_io_out_0_bits_isvec),
    .io_out_0_bits_sel_alu3(ibuffer_io_out_0_bits_sel_alu3),
    .io_out_0_bits_mask(ibuffer_io_out_0_bits_mask),
    .io_out_0_bits_sel_imm(ibuffer_io_out_0_bits_sel_imm),
    .io_out_0_bits_mem_unsigned(ibuffer_io_out_0_bits_mem_unsigned),
    .io_out_0_bits_alu_fn(ibuffer_io_out_0_bits_alu_fn),
    .io_out_0_bits_mem(ibuffer_io_out_0_bits_mem),
    .io_out_0_bits_mem_cmd(ibuffer_io_out_0_bits_mem_cmd),
    .io_out_0_bits_mop(ibuffer_io_out_0_bits_mop),
    .io_out_0_bits_reg_idx1(ibuffer_io_out_0_bits_reg_idx1),
    .io_out_0_bits_reg_idx2(ibuffer_io_out_0_bits_reg_idx2),
    .io_out_0_bits_reg_idx3(ibuffer_io_out_0_bits_reg_idx3),
    .io_out_0_bits_reg_idxw(ibuffer_io_out_0_bits_reg_idxw),
    .io_out_0_bits_wfd(ibuffer_io_out_0_bits_wfd),
    .io_out_0_bits_fence(ibuffer_io_out_0_bits_fence),
    .io_out_0_bits_sfu(ibuffer_io_out_0_bits_sfu),
    .io_out_0_bits_readmask(ibuffer_io_out_0_bits_readmask),
    .io_out_0_bits_writemask(ibuffer_io_out_0_bits_writemask),
    .io_out_0_bits_wxd(ibuffer_io_out_0_bits_wxd),
    .io_out_0_bits_pc(ibuffer_io_out_0_bits_pc),
    .io_out_1_ready(ibuffer_io_out_1_ready),
    .io_out_1_valid(ibuffer_io_out_1_valid),
    .io_out_1_bits_inst(ibuffer_io_out_1_bits_inst),
    .io_out_1_bits_wid(ibuffer_io_out_1_bits_wid),
    .io_out_1_bits_fp(ibuffer_io_out_1_bits_fp),
    .io_out_1_bits_branch(ibuffer_io_out_1_bits_branch),
    .io_out_1_bits_simt_stack(ibuffer_io_out_1_bits_simt_stack),
    .io_out_1_bits_simt_stack_op(ibuffer_io_out_1_bits_simt_stack_op),
    .io_out_1_bits_barrier(ibuffer_io_out_1_bits_barrier),
    .io_out_1_bits_csr(ibuffer_io_out_1_bits_csr),
    .io_out_1_bits_reverse(ibuffer_io_out_1_bits_reverse),
    .io_out_1_bits_sel_alu2(ibuffer_io_out_1_bits_sel_alu2),
    .io_out_1_bits_sel_alu1(ibuffer_io_out_1_bits_sel_alu1),
    .io_out_1_bits_isvec(ibuffer_io_out_1_bits_isvec),
    .io_out_1_bits_sel_alu3(ibuffer_io_out_1_bits_sel_alu3),
    .io_out_1_bits_mask(ibuffer_io_out_1_bits_mask),
    .io_out_1_bits_sel_imm(ibuffer_io_out_1_bits_sel_imm),
    .io_out_1_bits_mem_unsigned(ibuffer_io_out_1_bits_mem_unsigned),
    .io_out_1_bits_alu_fn(ibuffer_io_out_1_bits_alu_fn),
    .io_out_1_bits_mem(ibuffer_io_out_1_bits_mem),
    .io_out_1_bits_mem_cmd(ibuffer_io_out_1_bits_mem_cmd),
    .io_out_1_bits_mop(ibuffer_io_out_1_bits_mop),
    .io_out_1_bits_reg_idx1(ibuffer_io_out_1_bits_reg_idx1),
    .io_out_1_bits_reg_idx2(ibuffer_io_out_1_bits_reg_idx2),
    .io_out_1_bits_reg_idx3(ibuffer_io_out_1_bits_reg_idx3),
    .io_out_1_bits_reg_idxw(ibuffer_io_out_1_bits_reg_idxw),
    .io_out_1_bits_wfd(ibuffer_io_out_1_bits_wfd),
    .io_out_1_bits_fence(ibuffer_io_out_1_bits_fence),
    .io_out_1_bits_sfu(ibuffer_io_out_1_bits_sfu),
    .io_out_1_bits_readmask(ibuffer_io_out_1_bits_readmask),
    .io_out_1_bits_writemask(ibuffer_io_out_1_bits_writemask),
    .io_out_1_bits_wxd(ibuffer_io_out_1_bits_wxd),
    .io_out_1_bits_pc(ibuffer_io_out_1_bits_pc),
    .io_out_2_ready(ibuffer_io_out_2_ready),
    .io_out_2_valid(ibuffer_io_out_2_valid),
    .io_out_2_bits_inst(ibuffer_io_out_2_bits_inst),
    .io_out_2_bits_wid(ibuffer_io_out_2_bits_wid),
    .io_out_2_bits_fp(ibuffer_io_out_2_bits_fp),
    .io_out_2_bits_branch(ibuffer_io_out_2_bits_branch),
    .io_out_2_bits_simt_stack(ibuffer_io_out_2_bits_simt_stack),
    .io_out_2_bits_simt_stack_op(ibuffer_io_out_2_bits_simt_stack_op),
    .io_out_2_bits_barrier(ibuffer_io_out_2_bits_barrier),
    .io_out_2_bits_csr(ibuffer_io_out_2_bits_csr),
    .io_out_2_bits_reverse(ibuffer_io_out_2_bits_reverse),
    .io_out_2_bits_sel_alu2(ibuffer_io_out_2_bits_sel_alu2),
    .io_out_2_bits_sel_alu1(ibuffer_io_out_2_bits_sel_alu1),
    .io_out_2_bits_isvec(ibuffer_io_out_2_bits_isvec),
    .io_out_2_bits_sel_alu3(ibuffer_io_out_2_bits_sel_alu3),
    .io_out_2_bits_mask(ibuffer_io_out_2_bits_mask),
    .io_out_2_bits_sel_imm(ibuffer_io_out_2_bits_sel_imm),
    .io_out_2_bits_mem_unsigned(ibuffer_io_out_2_bits_mem_unsigned),
    .io_out_2_bits_alu_fn(ibuffer_io_out_2_bits_alu_fn),
    .io_out_2_bits_mem(ibuffer_io_out_2_bits_mem),
    .io_out_2_bits_mem_cmd(ibuffer_io_out_2_bits_mem_cmd),
    .io_out_2_bits_mop(ibuffer_io_out_2_bits_mop),
    .io_out_2_bits_reg_idx1(ibuffer_io_out_2_bits_reg_idx1),
    .io_out_2_bits_reg_idx2(ibuffer_io_out_2_bits_reg_idx2),
    .io_out_2_bits_reg_idx3(ibuffer_io_out_2_bits_reg_idx3),
    .io_out_2_bits_reg_idxw(ibuffer_io_out_2_bits_reg_idxw),
    .io_out_2_bits_wfd(ibuffer_io_out_2_bits_wfd),
    .io_out_2_bits_fence(ibuffer_io_out_2_bits_fence),
    .io_out_2_bits_sfu(ibuffer_io_out_2_bits_sfu),
    .io_out_2_bits_readmask(ibuffer_io_out_2_bits_readmask),
    .io_out_2_bits_writemask(ibuffer_io_out_2_bits_writemask),
    .io_out_2_bits_wxd(ibuffer_io_out_2_bits_wxd),
    .io_out_2_bits_pc(ibuffer_io_out_2_bits_pc),
    .io_out_3_ready(ibuffer_io_out_3_ready),
    .io_out_3_valid(ibuffer_io_out_3_valid),
    .io_out_3_bits_inst(ibuffer_io_out_3_bits_inst),
    .io_out_3_bits_wid(ibuffer_io_out_3_bits_wid),
    .io_out_3_bits_fp(ibuffer_io_out_3_bits_fp),
    .io_out_3_bits_branch(ibuffer_io_out_3_bits_branch),
    .io_out_3_bits_simt_stack(ibuffer_io_out_3_bits_simt_stack),
    .io_out_3_bits_simt_stack_op(ibuffer_io_out_3_bits_simt_stack_op),
    .io_out_3_bits_barrier(ibuffer_io_out_3_bits_barrier),
    .io_out_3_bits_csr(ibuffer_io_out_3_bits_csr),
    .io_out_3_bits_reverse(ibuffer_io_out_3_bits_reverse),
    .io_out_3_bits_sel_alu2(ibuffer_io_out_3_bits_sel_alu2),
    .io_out_3_bits_sel_alu1(ibuffer_io_out_3_bits_sel_alu1),
    .io_out_3_bits_isvec(ibuffer_io_out_3_bits_isvec),
    .io_out_3_bits_sel_alu3(ibuffer_io_out_3_bits_sel_alu3),
    .io_out_3_bits_mask(ibuffer_io_out_3_bits_mask),
    .io_out_3_bits_sel_imm(ibuffer_io_out_3_bits_sel_imm),
    .io_out_3_bits_mem_unsigned(ibuffer_io_out_3_bits_mem_unsigned),
    .io_out_3_bits_alu_fn(ibuffer_io_out_3_bits_alu_fn),
    .io_out_3_bits_mem(ibuffer_io_out_3_bits_mem),
    .io_out_3_bits_mem_cmd(ibuffer_io_out_3_bits_mem_cmd),
    .io_out_3_bits_mop(ibuffer_io_out_3_bits_mop),
    .io_out_3_bits_reg_idx1(ibuffer_io_out_3_bits_reg_idx1),
    .io_out_3_bits_reg_idx2(ibuffer_io_out_3_bits_reg_idx2),
    .io_out_3_bits_reg_idx3(ibuffer_io_out_3_bits_reg_idx3),
    .io_out_3_bits_reg_idxw(ibuffer_io_out_3_bits_reg_idxw),
    .io_out_3_bits_wfd(ibuffer_io_out_3_bits_wfd),
    .io_out_3_bits_fence(ibuffer_io_out_3_bits_fence),
    .io_out_3_bits_sfu(ibuffer_io_out_3_bits_sfu),
    .io_out_3_bits_readmask(ibuffer_io_out_3_bits_readmask),
    .io_out_3_bits_writemask(ibuffer_io_out_3_bits_writemask),
    .io_out_3_bits_wxd(ibuffer_io_out_3_bits_wxd),
    .io_out_3_bits_pc(ibuffer_io_out_3_bits_pc),
    .io_ibuffer_ready_0(ibuffer_io_ibuffer_ready_0),
    .io_ibuffer_ready_1(ibuffer_io_ibuffer_ready_1),
    .io_ibuffer_ready_2(ibuffer_io_ibuffer_ready_2),
    .io_ibuffer_ready_3(ibuffer_io_ibuffer_ready_3)
  );
  ibuffer2issue ibuffer2issue ( // @[pipe.scala 54:27]
    .clock(ibuffer2issue_clock),
    .io_in_0_ready(ibuffer2issue_io_in_0_ready),
    .io_in_0_valid(ibuffer2issue_io_in_0_valid),
    .io_in_0_bits_inst(ibuffer2issue_io_in_0_bits_inst),
    .io_in_0_bits_wid(ibuffer2issue_io_in_0_bits_wid),
    .io_in_0_bits_fp(ibuffer2issue_io_in_0_bits_fp),
    .io_in_0_bits_branch(ibuffer2issue_io_in_0_bits_branch),
    .io_in_0_bits_simt_stack(ibuffer2issue_io_in_0_bits_simt_stack),
    .io_in_0_bits_simt_stack_op(ibuffer2issue_io_in_0_bits_simt_stack_op),
    .io_in_0_bits_barrier(ibuffer2issue_io_in_0_bits_barrier),
    .io_in_0_bits_csr(ibuffer2issue_io_in_0_bits_csr),
    .io_in_0_bits_reverse(ibuffer2issue_io_in_0_bits_reverse),
    .io_in_0_bits_sel_alu2(ibuffer2issue_io_in_0_bits_sel_alu2),
    .io_in_0_bits_sel_alu1(ibuffer2issue_io_in_0_bits_sel_alu1),
    .io_in_0_bits_isvec(ibuffer2issue_io_in_0_bits_isvec),
    .io_in_0_bits_sel_alu3(ibuffer2issue_io_in_0_bits_sel_alu3),
    .io_in_0_bits_mask(ibuffer2issue_io_in_0_bits_mask),
    .io_in_0_bits_sel_imm(ibuffer2issue_io_in_0_bits_sel_imm),
    .io_in_0_bits_mem_unsigned(ibuffer2issue_io_in_0_bits_mem_unsigned),
    .io_in_0_bits_alu_fn(ibuffer2issue_io_in_0_bits_alu_fn),
    .io_in_0_bits_mem(ibuffer2issue_io_in_0_bits_mem),
    .io_in_0_bits_mem_cmd(ibuffer2issue_io_in_0_bits_mem_cmd),
    .io_in_0_bits_mop(ibuffer2issue_io_in_0_bits_mop),
    .io_in_0_bits_reg_idx1(ibuffer2issue_io_in_0_bits_reg_idx1),
    .io_in_0_bits_reg_idx2(ibuffer2issue_io_in_0_bits_reg_idx2),
    .io_in_0_bits_reg_idx3(ibuffer2issue_io_in_0_bits_reg_idx3),
    .io_in_0_bits_reg_idxw(ibuffer2issue_io_in_0_bits_reg_idxw),
    .io_in_0_bits_wfd(ibuffer2issue_io_in_0_bits_wfd),
    .io_in_0_bits_fence(ibuffer2issue_io_in_0_bits_fence),
    .io_in_0_bits_sfu(ibuffer2issue_io_in_0_bits_sfu),
    .io_in_0_bits_readmask(ibuffer2issue_io_in_0_bits_readmask),
    .io_in_0_bits_writemask(ibuffer2issue_io_in_0_bits_writemask),
    .io_in_0_bits_wxd(ibuffer2issue_io_in_0_bits_wxd),
    .io_in_0_bits_pc(ibuffer2issue_io_in_0_bits_pc),
    .io_in_1_ready(ibuffer2issue_io_in_1_ready),
    .io_in_1_valid(ibuffer2issue_io_in_1_valid),
    .io_in_1_bits_inst(ibuffer2issue_io_in_1_bits_inst),
    .io_in_1_bits_wid(ibuffer2issue_io_in_1_bits_wid),
    .io_in_1_bits_fp(ibuffer2issue_io_in_1_bits_fp),
    .io_in_1_bits_branch(ibuffer2issue_io_in_1_bits_branch),
    .io_in_1_bits_simt_stack(ibuffer2issue_io_in_1_bits_simt_stack),
    .io_in_1_bits_simt_stack_op(ibuffer2issue_io_in_1_bits_simt_stack_op),
    .io_in_1_bits_barrier(ibuffer2issue_io_in_1_bits_barrier),
    .io_in_1_bits_csr(ibuffer2issue_io_in_1_bits_csr),
    .io_in_1_bits_reverse(ibuffer2issue_io_in_1_bits_reverse),
    .io_in_1_bits_sel_alu2(ibuffer2issue_io_in_1_bits_sel_alu2),
    .io_in_1_bits_sel_alu1(ibuffer2issue_io_in_1_bits_sel_alu1),
    .io_in_1_bits_isvec(ibuffer2issue_io_in_1_bits_isvec),
    .io_in_1_bits_sel_alu3(ibuffer2issue_io_in_1_bits_sel_alu3),
    .io_in_1_bits_mask(ibuffer2issue_io_in_1_bits_mask),
    .io_in_1_bits_sel_imm(ibuffer2issue_io_in_1_bits_sel_imm),
    .io_in_1_bits_mem_unsigned(ibuffer2issue_io_in_1_bits_mem_unsigned),
    .io_in_1_bits_alu_fn(ibuffer2issue_io_in_1_bits_alu_fn),
    .io_in_1_bits_mem(ibuffer2issue_io_in_1_bits_mem),
    .io_in_1_bits_mem_cmd(ibuffer2issue_io_in_1_bits_mem_cmd),
    .io_in_1_bits_mop(ibuffer2issue_io_in_1_bits_mop),
    .io_in_1_bits_reg_idx1(ibuffer2issue_io_in_1_bits_reg_idx1),
    .io_in_1_bits_reg_idx2(ibuffer2issue_io_in_1_bits_reg_idx2),
    .io_in_1_bits_reg_idx3(ibuffer2issue_io_in_1_bits_reg_idx3),
    .io_in_1_bits_reg_idxw(ibuffer2issue_io_in_1_bits_reg_idxw),
    .io_in_1_bits_wfd(ibuffer2issue_io_in_1_bits_wfd),
    .io_in_1_bits_fence(ibuffer2issue_io_in_1_bits_fence),
    .io_in_1_bits_sfu(ibuffer2issue_io_in_1_bits_sfu),
    .io_in_1_bits_readmask(ibuffer2issue_io_in_1_bits_readmask),
    .io_in_1_bits_writemask(ibuffer2issue_io_in_1_bits_writemask),
    .io_in_1_bits_wxd(ibuffer2issue_io_in_1_bits_wxd),
    .io_in_1_bits_pc(ibuffer2issue_io_in_1_bits_pc),
    .io_in_2_ready(ibuffer2issue_io_in_2_ready),
    .io_in_2_valid(ibuffer2issue_io_in_2_valid),
    .io_in_2_bits_inst(ibuffer2issue_io_in_2_bits_inst),
    .io_in_2_bits_wid(ibuffer2issue_io_in_2_bits_wid),
    .io_in_2_bits_fp(ibuffer2issue_io_in_2_bits_fp),
    .io_in_2_bits_branch(ibuffer2issue_io_in_2_bits_branch),
    .io_in_2_bits_simt_stack(ibuffer2issue_io_in_2_bits_simt_stack),
    .io_in_2_bits_simt_stack_op(ibuffer2issue_io_in_2_bits_simt_stack_op),
    .io_in_2_bits_barrier(ibuffer2issue_io_in_2_bits_barrier),
    .io_in_2_bits_csr(ibuffer2issue_io_in_2_bits_csr),
    .io_in_2_bits_reverse(ibuffer2issue_io_in_2_bits_reverse),
    .io_in_2_bits_sel_alu2(ibuffer2issue_io_in_2_bits_sel_alu2),
    .io_in_2_bits_sel_alu1(ibuffer2issue_io_in_2_bits_sel_alu1),
    .io_in_2_bits_isvec(ibuffer2issue_io_in_2_bits_isvec),
    .io_in_2_bits_sel_alu3(ibuffer2issue_io_in_2_bits_sel_alu3),
    .io_in_2_bits_mask(ibuffer2issue_io_in_2_bits_mask),
    .io_in_2_bits_sel_imm(ibuffer2issue_io_in_2_bits_sel_imm),
    .io_in_2_bits_mem_unsigned(ibuffer2issue_io_in_2_bits_mem_unsigned),
    .io_in_2_bits_alu_fn(ibuffer2issue_io_in_2_bits_alu_fn),
    .io_in_2_bits_mem(ibuffer2issue_io_in_2_bits_mem),
    .io_in_2_bits_mem_cmd(ibuffer2issue_io_in_2_bits_mem_cmd),
    .io_in_2_bits_mop(ibuffer2issue_io_in_2_bits_mop),
    .io_in_2_bits_reg_idx1(ibuffer2issue_io_in_2_bits_reg_idx1),
    .io_in_2_bits_reg_idx2(ibuffer2issue_io_in_2_bits_reg_idx2),
    .io_in_2_bits_reg_idx3(ibuffer2issue_io_in_2_bits_reg_idx3),
    .io_in_2_bits_reg_idxw(ibuffer2issue_io_in_2_bits_reg_idxw),
    .io_in_2_bits_wfd(ibuffer2issue_io_in_2_bits_wfd),
    .io_in_2_bits_fence(ibuffer2issue_io_in_2_bits_fence),
    .io_in_2_bits_sfu(ibuffer2issue_io_in_2_bits_sfu),
    .io_in_2_bits_readmask(ibuffer2issue_io_in_2_bits_readmask),
    .io_in_2_bits_writemask(ibuffer2issue_io_in_2_bits_writemask),
    .io_in_2_bits_wxd(ibuffer2issue_io_in_2_bits_wxd),
    .io_in_2_bits_pc(ibuffer2issue_io_in_2_bits_pc),
    .io_in_3_ready(ibuffer2issue_io_in_3_ready),
    .io_in_3_valid(ibuffer2issue_io_in_3_valid),
    .io_in_3_bits_inst(ibuffer2issue_io_in_3_bits_inst),
    .io_in_3_bits_wid(ibuffer2issue_io_in_3_bits_wid),
    .io_in_3_bits_fp(ibuffer2issue_io_in_3_bits_fp),
    .io_in_3_bits_branch(ibuffer2issue_io_in_3_bits_branch),
    .io_in_3_bits_simt_stack(ibuffer2issue_io_in_3_bits_simt_stack),
    .io_in_3_bits_simt_stack_op(ibuffer2issue_io_in_3_bits_simt_stack_op),
    .io_in_3_bits_barrier(ibuffer2issue_io_in_3_bits_barrier),
    .io_in_3_bits_csr(ibuffer2issue_io_in_3_bits_csr),
    .io_in_3_bits_reverse(ibuffer2issue_io_in_3_bits_reverse),
    .io_in_3_bits_sel_alu2(ibuffer2issue_io_in_3_bits_sel_alu2),
    .io_in_3_bits_sel_alu1(ibuffer2issue_io_in_3_bits_sel_alu1),
    .io_in_3_bits_isvec(ibuffer2issue_io_in_3_bits_isvec),
    .io_in_3_bits_sel_alu3(ibuffer2issue_io_in_3_bits_sel_alu3),
    .io_in_3_bits_mask(ibuffer2issue_io_in_3_bits_mask),
    .io_in_3_bits_sel_imm(ibuffer2issue_io_in_3_bits_sel_imm),
    .io_in_3_bits_mem_unsigned(ibuffer2issue_io_in_3_bits_mem_unsigned),
    .io_in_3_bits_alu_fn(ibuffer2issue_io_in_3_bits_alu_fn),
    .io_in_3_bits_mem(ibuffer2issue_io_in_3_bits_mem),
    .io_in_3_bits_mem_cmd(ibuffer2issue_io_in_3_bits_mem_cmd),
    .io_in_3_bits_mop(ibuffer2issue_io_in_3_bits_mop),
    .io_in_3_bits_reg_idx1(ibuffer2issue_io_in_3_bits_reg_idx1),
    .io_in_3_bits_reg_idx2(ibuffer2issue_io_in_3_bits_reg_idx2),
    .io_in_3_bits_reg_idx3(ibuffer2issue_io_in_3_bits_reg_idx3),
    .io_in_3_bits_reg_idxw(ibuffer2issue_io_in_3_bits_reg_idxw),
    .io_in_3_bits_wfd(ibuffer2issue_io_in_3_bits_wfd),
    .io_in_3_bits_fence(ibuffer2issue_io_in_3_bits_fence),
    .io_in_3_bits_sfu(ibuffer2issue_io_in_3_bits_sfu),
    .io_in_3_bits_readmask(ibuffer2issue_io_in_3_bits_readmask),
    .io_in_3_bits_writemask(ibuffer2issue_io_in_3_bits_writemask),
    .io_in_3_bits_wxd(ibuffer2issue_io_in_3_bits_wxd),
    .io_in_3_bits_pc(ibuffer2issue_io_in_3_bits_pc),
    .io_out_ready(ibuffer2issue_io_out_ready),
    .io_out_valid(ibuffer2issue_io_out_valid),
    .io_out_bits_inst(ibuffer2issue_io_out_bits_inst),
    .io_out_bits_wid(ibuffer2issue_io_out_bits_wid),
    .io_out_bits_fp(ibuffer2issue_io_out_bits_fp),
    .io_out_bits_branch(ibuffer2issue_io_out_bits_branch),
    .io_out_bits_simt_stack(ibuffer2issue_io_out_bits_simt_stack),
    .io_out_bits_simt_stack_op(ibuffer2issue_io_out_bits_simt_stack_op),
    .io_out_bits_barrier(ibuffer2issue_io_out_bits_barrier),
    .io_out_bits_csr(ibuffer2issue_io_out_bits_csr),
    .io_out_bits_reverse(ibuffer2issue_io_out_bits_reverse),
    .io_out_bits_sel_alu2(ibuffer2issue_io_out_bits_sel_alu2),
    .io_out_bits_sel_alu1(ibuffer2issue_io_out_bits_sel_alu1),
    .io_out_bits_isvec(ibuffer2issue_io_out_bits_isvec),
    .io_out_bits_sel_alu3(ibuffer2issue_io_out_bits_sel_alu3),
    .io_out_bits_mask(ibuffer2issue_io_out_bits_mask),
    .io_out_bits_sel_imm(ibuffer2issue_io_out_bits_sel_imm),
    .io_out_bits_mem_unsigned(ibuffer2issue_io_out_bits_mem_unsigned),
    .io_out_bits_alu_fn(ibuffer2issue_io_out_bits_alu_fn),
    .io_out_bits_mem(ibuffer2issue_io_out_bits_mem),
    .io_out_bits_mem_cmd(ibuffer2issue_io_out_bits_mem_cmd),
    .io_out_bits_mop(ibuffer2issue_io_out_bits_mop),
    .io_out_bits_reg_idx1(ibuffer2issue_io_out_bits_reg_idx1),
    .io_out_bits_reg_idx2(ibuffer2issue_io_out_bits_reg_idx2),
    .io_out_bits_reg_idx3(ibuffer2issue_io_out_bits_reg_idx3),
    .io_out_bits_reg_idxw(ibuffer2issue_io_out_bits_reg_idxw),
    .io_out_bits_wfd(ibuffer2issue_io_out_bits_wfd),
    .io_out_bits_fence(ibuffer2issue_io_out_bits_fence),
    .io_out_bits_sfu(ibuffer2issue_io_out_bits_sfu),
    .io_out_bits_readmask(ibuffer2issue_io_out_bits_readmask),
    .io_out_bits_writemask(ibuffer2issue_io_out_bits_writemask),
    .io_out_bits_wxd(ibuffer2issue_io_out_bits_wxd),
    .io_out_bits_pc(ibuffer2issue_io_out_bits_pc)
  );
  Queue_41 exe_data ( // @[pipe.scala 55:22]
    .clock(exe_data_clock),
    .reset(exe_data_reset),
    .io_enq_ready(exe_data_io_enq_ready),
    .io_enq_valid(exe_data_io_enq_valid),
    .io_enq_bits_in1_0(exe_data_io_enq_bits_in1_0),
    .io_enq_bits_in1_1(exe_data_io_enq_bits_in1_1),
    .io_enq_bits_in1_2(exe_data_io_enq_bits_in1_2),
    .io_enq_bits_in1_3(exe_data_io_enq_bits_in1_3),
    .io_enq_bits_in1_4(exe_data_io_enq_bits_in1_4),
    .io_enq_bits_in1_5(exe_data_io_enq_bits_in1_5),
    .io_enq_bits_in1_6(exe_data_io_enq_bits_in1_6),
    .io_enq_bits_in1_7(exe_data_io_enq_bits_in1_7),
    .io_enq_bits_in2_0(exe_data_io_enq_bits_in2_0),
    .io_enq_bits_in2_1(exe_data_io_enq_bits_in2_1),
    .io_enq_bits_in2_2(exe_data_io_enq_bits_in2_2),
    .io_enq_bits_in2_3(exe_data_io_enq_bits_in2_3),
    .io_enq_bits_in2_4(exe_data_io_enq_bits_in2_4),
    .io_enq_bits_in2_5(exe_data_io_enq_bits_in2_5),
    .io_enq_bits_in2_6(exe_data_io_enq_bits_in2_6),
    .io_enq_bits_in2_7(exe_data_io_enq_bits_in2_7),
    .io_enq_bits_in3_0(exe_data_io_enq_bits_in3_0),
    .io_enq_bits_in3_1(exe_data_io_enq_bits_in3_1),
    .io_enq_bits_in3_2(exe_data_io_enq_bits_in3_2),
    .io_enq_bits_in3_3(exe_data_io_enq_bits_in3_3),
    .io_enq_bits_in3_4(exe_data_io_enq_bits_in3_4),
    .io_enq_bits_in3_5(exe_data_io_enq_bits_in3_5),
    .io_enq_bits_in3_6(exe_data_io_enq_bits_in3_6),
    .io_enq_bits_in3_7(exe_data_io_enq_bits_in3_7),
    .io_enq_bits_mask_0(exe_data_io_enq_bits_mask_0),
    .io_enq_bits_mask_1(exe_data_io_enq_bits_mask_1),
    .io_enq_bits_mask_2(exe_data_io_enq_bits_mask_2),
    .io_enq_bits_mask_3(exe_data_io_enq_bits_mask_3),
    .io_enq_bits_mask_4(exe_data_io_enq_bits_mask_4),
    .io_enq_bits_mask_5(exe_data_io_enq_bits_mask_5),
    .io_enq_bits_mask_6(exe_data_io_enq_bits_mask_6),
    .io_enq_bits_mask_7(exe_data_io_enq_bits_mask_7),
    .io_enq_bits_ctrl_inst(exe_data_io_enq_bits_ctrl_inst),
    .io_enq_bits_ctrl_wid(exe_data_io_enq_bits_ctrl_wid),
    .io_enq_bits_ctrl_fp(exe_data_io_enq_bits_ctrl_fp),
    .io_enq_bits_ctrl_branch(exe_data_io_enq_bits_ctrl_branch),
    .io_enq_bits_ctrl_simt_stack(exe_data_io_enq_bits_ctrl_simt_stack),
    .io_enq_bits_ctrl_simt_stack_op(exe_data_io_enq_bits_ctrl_simt_stack_op),
    .io_enq_bits_ctrl_barrier(exe_data_io_enq_bits_ctrl_barrier),
    .io_enq_bits_ctrl_csr(exe_data_io_enq_bits_ctrl_csr),
    .io_enq_bits_ctrl_reverse(exe_data_io_enq_bits_ctrl_reverse),
    .io_enq_bits_ctrl_isvec(exe_data_io_enq_bits_ctrl_isvec),
    .io_enq_bits_ctrl_mem_unsigned(exe_data_io_enq_bits_ctrl_mem_unsigned),
    .io_enq_bits_ctrl_alu_fn(exe_data_io_enq_bits_ctrl_alu_fn),
    .io_enq_bits_ctrl_mem(exe_data_io_enq_bits_ctrl_mem),
    .io_enq_bits_ctrl_mem_cmd(exe_data_io_enq_bits_ctrl_mem_cmd),
    .io_enq_bits_ctrl_mop(exe_data_io_enq_bits_ctrl_mop),
    .io_enq_bits_ctrl_reg_idxw(exe_data_io_enq_bits_ctrl_reg_idxw),
    .io_enq_bits_ctrl_wfd(exe_data_io_enq_bits_ctrl_wfd),
    .io_enq_bits_ctrl_fence(exe_data_io_enq_bits_ctrl_fence),
    .io_enq_bits_ctrl_sfu(exe_data_io_enq_bits_ctrl_sfu),
    .io_enq_bits_ctrl_readmask(exe_data_io_enq_bits_ctrl_readmask),
    .io_enq_bits_ctrl_writemask(exe_data_io_enq_bits_ctrl_writemask),
    .io_enq_bits_ctrl_wxd(exe_data_io_enq_bits_ctrl_wxd),
    .io_enq_bits_ctrl_pc(exe_data_io_enq_bits_ctrl_pc),
    .io_deq_ready(exe_data_io_deq_ready),
    .io_deq_valid(exe_data_io_deq_valid),
    .io_deq_bits_in1_0(exe_data_io_deq_bits_in1_0),
    .io_deq_bits_in1_1(exe_data_io_deq_bits_in1_1),
    .io_deq_bits_in1_2(exe_data_io_deq_bits_in1_2),
    .io_deq_bits_in1_3(exe_data_io_deq_bits_in1_3),
    .io_deq_bits_in1_4(exe_data_io_deq_bits_in1_4),
    .io_deq_bits_in1_5(exe_data_io_deq_bits_in1_5),
    .io_deq_bits_in1_6(exe_data_io_deq_bits_in1_6),
    .io_deq_bits_in1_7(exe_data_io_deq_bits_in1_7),
    .io_deq_bits_in2_0(exe_data_io_deq_bits_in2_0),
    .io_deq_bits_in2_1(exe_data_io_deq_bits_in2_1),
    .io_deq_bits_in2_2(exe_data_io_deq_bits_in2_2),
    .io_deq_bits_in2_3(exe_data_io_deq_bits_in2_3),
    .io_deq_bits_in2_4(exe_data_io_deq_bits_in2_4),
    .io_deq_bits_in2_5(exe_data_io_deq_bits_in2_5),
    .io_deq_bits_in2_6(exe_data_io_deq_bits_in2_6),
    .io_deq_bits_in2_7(exe_data_io_deq_bits_in2_7),
    .io_deq_bits_in3_0(exe_data_io_deq_bits_in3_0),
    .io_deq_bits_in3_1(exe_data_io_deq_bits_in3_1),
    .io_deq_bits_in3_2(exe_data_io_deq_bits_in3_2),
    .io_deq_bits_in3_3(exe_data_io_deq_bits_in3_3),
    .io_deq_bits_in3_4(exe_data_io_deq_bits_in3_4),
    .io_deq_bits_in3_5(exe_data_io_deq_bits_in3_5),
    .io_deq_bits_in3_6(exe_data_io_deq_bits_in3_6),
    .io_deq_bits_in3_7(exe_data_io_deq_bits_in3_7),
    .io_deq_bits_mask_0(exe_data_io_deq_bits_mask_0),
    .io_deq_bits_mask_1(exe_data_io_deq_bits_mask_1),
    .io_deq_bits_mask_2(exe_data_io_deq_bits_mask_2),
    .io_deq_bits_mask_3(exe_data_io_deq_bits_mask_3),
    .io_deq_bits_mask_4(exe_data_io_deq_bits_mask_4),
    .io_deq_bits_mask_5(exe_data_io_deq_bits_mask_5),
    .io_deq_bits_mask_6(exe_data_io_deq_bits_mask_6),
    .io_deq_bits_mask_7(exe_data_io_deq_bits_mask_7),
    .io_deq_bits_ctrl_inst(exe_data_io_deq_bits_ctrl_inst),
    .io_deq_bits_ctrl_wid(exe_data_io_deq_bits_ctrl_wid),
    .io_deq_bits_ctrl_fp(exe_data_io_deq_bits_ctrl_fp),
    .io_deq_bits_ctrl_branch(exe_data_io_deq_bits_ctrl_branch),
    .io_deq_bits_ctrl_simt_stack(exe_data_io_deq_bits_ctrl_simt_stack),
    .io_deq_bits_ctrl_simt_stack_op(exe_data_io_deq_bits_ctrl_simt_stack_op),
    .io_deq_bits_ctrl_barrier(exe_data_io_deq_bits_ctrl_barrier),
    .io_deq_bits_ctrl_csr(exe_data_io_deq_bits_ctrl_csr),
    .io_deq_bits_ctrl_reverse(exe_data_io_deq_bits_ctrl_reverse),
    .io_deq_bits_ctrl_isvec(exe_data_io_deq_bits_ctrl_isvec),
    .io_deq_bits_ctrl_mem_unsigned(exe_data_io_deq_bits_ctrl_mem_unsigned),
    .io_deq_bits_ctrl_alu_fn(exe_data_io_deq_bits_ctrl_alu_fn),
    .io_deq_bits_ctrl_mem(exe_data_io_deq_bits_ctrl_mem),
    .io_deq_bits_ctrl_mem_cmd(exe_data_io_deq_bits_ctrl_mem_cmd),
    .io_deq_bits_ctrl_mop(exe_data_io_deq_bits_ctrl_mop),
    .io_deq_bits_ctrl_reg_idxw(exe_data_io_deq_bits_ctrl_reg_idxw),
    .io_deq_bits_ctrl_wfd(exe_data_io_deq_bits_ctrl_wfd),
    .io_deq_bits_ctrl_fence(exe_data_io_deq_bits_ctrl_fence),
    .io_deq_bits_ctrl_sfu(exe_data_io_deq_bits_ctrl_sfu),
    .io_deq_bits_ctrl_readmask(exe_data_io_deq_bits_ctrl_readmask),
    .io_deq_bits_ctrl_writemask(exe_data_io_deq_bits_ctrl_writemask),
    .io_deq_bits_ctrl_wxd(exe_data_io_deq_bits_ctrl_wxd),
    .io_deq_bits_ctrl_pc(exe_data_io_deq_bits_ctrl_pc)
  );
  SIMT_STACK simt_stack ( // @[pipe.scala 56:24]
    .clock(simt_stack_clock),
    .reset(simt_stack_reset),
    .io_branch_ctl_ready(simt_stack_io_branch_ctl_ready),
    .io_branch_ctl_valid(simt_stack_io_branch_ctl_valid),
    .io_branch_ctl_bits_opcode(simt_stack_io_branch_ctl_bits_opcode),
    .io_branch_ctl_bits_wid(simt_stack_io_branch_ctl_bits_wid),
    .io_branch_ctl_bits_PC_branch(simt_stack_io_branch_ctl_bits_PC_branch),
    .io_branch_ctl_bits_mask_init(simt_stack_io_branch_ctl_bits_mask_init),
    .io_if_mask_ready(simt_stack_io_if_mask_ready),
    .io_if_mask_valid(simt_stack_io_if_mask_valid),
    .io_if_mask_bits_if_mask(simt_stack_io_if_mask_bits_if_mask),
    .io_if_mask_bits_wid(simt_stack_io_if_mask_bits_wid),
    .io_input_wid(simt_stack_io_input_wid),
    .io_out_mask(simt_stack_io_out_mask),
    .io_complete_valid(simt_stack_io_complete_valid),
    .io_complete_bits(simt_stack_io_complete_bits),
    .io_fetch_ctl_ready(simt_stack_io_fetch_ctl_ready),
    .io_fetch_ctl_valid(simt_stack_io_fetch_ctl_valid),
    .io_fetch_ctl_bits_wid(simt_stack_io_fetch_ctl_bits_wid),
    .io_fetch_ctl_bits_jump(simt_stack_io_fetch_ctl_bits_jump),
    .io_fetch_ctl_bits_new_pc(simt_stack_io_fetch_ctl_bits_new_pc)
  );
  Branch_back branch_back ( // @[pipe.scala 57:25]
    .io_out_ready(branch_back_io_out_ready),
    .io_out_valid(branch_back_io_out_valid),
    .io_out_bits_wid(branch_back_io_out_bits_wid),
    .io_out_bits_jump(branch_back_io_out_bits_jump),
    .io_out_bits_new_pc(branch_back_io_out_bits_new_pc),
    .io_in0_ready(branch_back_io_in0_ready),
    .io_in0_valid(branch_back_io_in0_valid),
    .io_in0_bits_wid(branch_back_io_in0_bits_wid),
    .io_in0_bits_jump(branch_back_io_in0_bits_jump),
    .io_in0_bits_new_pc(branch_back_io_in0_bits_new_pc),
    .io_in1_ready(branch_back_io_in1_ready),
    .io_in1_valid(branch_back_io_in1_valid),
    .io_in1_bits_wid(branch_back_io_in1_bits_wid),
    .io_in1_bits_jump(branch_back_io_in1_bits_jump),
    .io_in1_bits_new_pc(branch_back_io_in1_bits_new_pc)
  );
  CSRexe csrfile ( // @[pipe.scala 58:21]
    .clock(csrfile_clock),
    .reset(csrfile_reset),
    .io_in_ready(csrfile_io_in_ready),
    .io_in_valid(csrfile_io_in_valid),
    .io_in_bits_ctrl_inst(csrfile_io_in_bits_ctrl_inst),
    .io_in_bits_ctrl_wid(csrfile_io_in_bits_ctrl_wid),
    .io_in_bits_ctrl_csr(csrfile_io_in_bits_ctrl_csr),
    .io_in_bits_ctrl_isvec(csrfile_io_in_bits_ctrl_isvec),
    .io_in_bits_ctrl_reg_idxw(csrfile_io_in_bits_ctrl_reg_idxw),
    .io_in_bits_ctrl_wxd(csrfile_io_in_bits_ctrl_wxd),
    .io_in_bits_in1(csrfile_io_in_bits_in1),
    .io_out_ready(csrfile_io_out_ready),
    .io_out_valid(csrfile_io_out_valid),
    .io_out_bits_wb_wxd_rd(csrfile_io_out_bits_wb_wxd_rd),
    .io_out_bits_wxd(csrfile_io_out_bits_wxd),
    .io_out_bits_reg_idxw(csrfile_io_out_bits_reg_idxw),
    .io_out_bits_warp_id(csrfile_io_out_bits_warp_id),
    .io_frm_wid(csrfile_io_frm_wid),
    .io_frm(csrfile_io_frm),
    .io_CTA2csr_valid(csrfile_io_CTA2csr_valid),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count(csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch(csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch(csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch(csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch
      ),
    .io_CTA2csr_bits_wid(csrfile_io_CTA2csr_bits_wid)
  );
  assign io_icache_req_valid = warp_sche_io_pc_req_valid; // @[pipe.scala 73:22]
  assign io_icache_req_bits_addr = warp_sche_io_pc_req_bits_addr; // @[pipe.scala 73:22]
  assign io_icache_req_bits_warpid = warp_sche_io_pc_req_bits_warpid; // @[pipe.scala 73:22]
  assign io_externalFlushPipe_valid = warp_sche_io_flush_valid | warp_sche_io_flushCache_valid; // @[pipe.scala 60:55]
  assign io_externalFlushPipe_bits = warp_sche_io_flush_valid ? warp_sche_io_flush_bits : warp_sche_io_flushCache_bits; // @[pipe.scala 61:33]
  assign io_dcache_req_valid = lsu_io_dcache_req_valid; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_instrId = lsu_io_dcache_req_bits_instrId; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_isWrite = lsu_io_dcache_req_bits_isWrite; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_tag = lsu_io_dcache_req_bits_tag; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_setIdx = lsu_io_dcache_req_bits_setIdx; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_0_activeMask = lsu_io_dcache_req_bits_perLaneAddr_0_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_0_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_0_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_1_activeMask = lsu_io_dcache_req_bits_perLaneAddr_1_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_1_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_1_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_2_activeMask = lsu_io_dcache_req_bits_perLaneAddr_2_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_2_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_2_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_3_activeMask = lsu_io_dcache_req_bits_perLaneAddr_3_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_3_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_3_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_4_activeMask = lsu_io_dcache_req_bits_perLaneAddr_4_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_4_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_4_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_5_activeMask = lsu_io_dcache_req_bits_perLaneAddr_5_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_5_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_5_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_6_activeMask = lsu_io_dcache_req_bits_perLaneAddr_6_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_6_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_6_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_7_activeMask = lsu_io_dcache_req_bits_perLaneAddr_7_activeMask; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_perLaneAddr_7_blockOffset = lsu_io_dcache_req_bits_perLaneAddr_7_blockOffset; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_0 = lsu_io_dcache_req_bits_data_0; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_1 = lsu_io_dcache_req_bits_data_1; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_2 = lsu_io_dcache_req_bits_data_2; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_3 = lsu_io_dcache_req_bits_data_3; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_4 = lsu_io_dcache_req_bits_data_4; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_5 = lsu_io_dcache_req_bits_data_5; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_6 = lsu_io_dcache_req_bits_data_6; // @[pipe.scala 234:20]
  assign io_dcache_req_bits_data_7 = lsu_io_dcache_req_bits_data_7; // @[pipe.scala 234:20]
  assign io_dcache_rsp_ready = lsu_io_dcache_rsp_ready; // @[pipe.scala 233:20]
  assign io_shared_req_valid = lsu_io_shared_req_valid; // @[pipe.scala 237:20]
  assign io_shared_req_bits_instrId = lsu_io_shared_req_bits_instrId; // @[pipe.scala 237:20]
  assign io_shared_req_bits_isWrite = lsu_io_shared_req_bits_isWrite; // @[pipe.scala 237:20]
  assign io_shared_req_bits_setIdx = lsu_io_shared_req_bits_setIdx; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_0_activeMask = lsu_io_shared_req_bits_perLaneAddr_0_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_0_blockOffset = lsu_io_shared_req_bits_perLaneAddr_0_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_1_activeMask = lsu_io_shared_req_bits_perLaneAddr_1_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_1_blockOffset = lsu_io_shared_req_bits_perLaneAddr_1_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_2_activeMask = lsu_io_shared_req_bits_perLaneAddr_2_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_2_blockOffset = lsu_io_shared_req_bits_perLaneAddr_2_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_3_activeMask = lsu_io_shared_req_bits_perLaneAddr_3_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_3_blockOffset = lsu_io_shared_req_bits_perLaneAddr_3_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_4_activeMask = lsu_io_shared_req_bits_perLaneAddr_4_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_4_blockOffset = lsu_io_shared_req_bits_perLaneAddr_4_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_5_activeMask = lsu_io_shared_req_bits_perLaneAddr_5_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_5_blockOffset = lsu_io_shared_req_bits_perLaneAddr_5_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_6_activeMask = lsu_io_shared_req_bits_perLaneAddr_6_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_6_blockOffset = lsu_io_shared_req_bits_perLaneAddr_6_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_7_activeMask = lsu_io_shared_req_bits_perLaneAddr_7_activeMask; // @[pipe.scala 237:20]
  assign io_shared_req_bits_perLaneAddr_7_blockOffset = lsu_io_shared_req_bits_perLaneAddr_7_blockOffset; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_0 = lsu_io_shared_req_bits_data_0; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_1 = lsu_io_shared_req_bits_data_1; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_2 = lsu_io_shared_req_bits_data_2; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_3 = lsu_io_shared_req_bits_data_3; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_4 = lsu_io_shared_req_bits_data_4; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_5 = lsu_io_shared_req_bits_data_5; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_6 = lsu_io_shared_req_bits_data_6; // @[pipe.scala 237:20]
  assign io_shared_req_bits_data_7 = lsu_io_shared_req_bits_data_7; // @[pipe.scala 237:20]
  assign io_shared_rsp_ready = lsu_io_shared_rsp_ready; // @[pipe.scala 236:20]
  assign io_warpRsp_valid = warp_sche_io_warpRsp_valid; // @[pipe.scala 81:23]
  assign io_warpRsp_bits_wid = warp_sche_io_warpRsp_bits_wid; // @[pipe.scala 81:23]
  assign io_wg_id_lookup = warp_sche_io_wg_id_lookup; // @[pipe.scala 68:18]
  assign warp_sche_clock = clock;
  assign warp_sche_reset = reset;
  assign warp_sche_io_pc_reset = io_pc_reset; // @[pipe.scala 63:24]
  assign warp_sche_io_warpReq_valid = io_warpReq_valid; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count = io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch =
    io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch; // @[pipe.scala 80:23]
  assign warp_sche_io_warpReq_bits_wid = io_warpReq_bits_wid; // @[pipe.scala 80:23]
  assign warp_sche_io_wg_id_tag = io_wg_id_tag; // @[pipe.scala 67:25]
  assign warp_sche_io_pc_rsp_valid = io_icache_rsp_valid; // @[pipe.scala 69:28]
  assign warp_sche_io_pc_rsp_bits_addr = io_icache_rsp_bits_addr; // @[pipe.scala 70:27]
  assign warp_sche_io_pc_rsp_bits_warpid = io_icache_rsp_bits_warpid; // @[pipe.scala 70:27]
  assign warp_sche_io_pc_rsp_bits_status = ibuffer_io_in_ready ? io_icache_rsp_bits_status : 2'h1; // @[pipe.scala 71:39]
  assign warp_sche_io_branch_valid = branch_back_io_out_valid; // @[pipe.scala 64:22]
  assign warp_sche_io_branch_bits_wid = branch_back_io_out_bits_wid; // @[pipe.scala 64:22]
  assign warp_sche_io_branch_bits_jump = branch_back_io_out_bits_jump; // @[pipe.scala 64:22]
  assign warp_sche_io_branch_bits_new_pc = branch_back_io_out_bits_new_pc; // @[pipe.scala 64:22]
  assign warp_sche_io_warp_control_valid = issue_io_out_warpscheduler_valid; // @[pipe.scala 74:28]
  assign warp_sche_io_warp_control_bits_ctrl_wid = issue_io_out_warpscheduler_bits_ctrl_wid; // @[pipe.scala 74:28]
  assign warp_sche_io_warp_control_bits_ctrl_simt_stack_op = issue_io_out_warpscheduler_bits_ctrl_simt_stack_op; // @[pipe.scala 74:28]
  assign warp_sche_io_warp_control_bits_ctrl_barrier = issue_io_out_warpscheduler_bits_ctrl_barrier; // @[pipe.scala 74:28]
  assign warp_sche_io_scoreboard_busy = {warp_sche_io_scoreboard_busy_hi,warp_sche_io_scoreboard_busy_lo}; // @[pipe.scala 77:70]
  assign warp_sche_io_exe_busy = ~_warp_sche_io_exe_busy_T; // @[pipe.scala 116:27]
  assign warp_sche_io_pc_ibuffer_ready_0 = ibuffer_io_ibuffer_ready_0; // @[pipe.scala 66:32]
  assign warp_sche_io_pc_ibuffer_ready_1 = ibuffer_io_ibuffer_ready_1; // @[pipe.scala 66:32]
  assign warp_sche_io_pc_ibuffer_ready_2 = ibuffer_io_ibuffer_ready_2; // @[pipe.scala 66:32]
  assign warp_sche_io_pc_ibuffer_ready_3 = ibuffer_io_ibuffer_ready_3; // @[pipe.scala 66:32]
  assign control_io_inst = io_icache_rsp_bits_data; // @[pipe.scala 94:18]
  assign control_io_pc = io_icache_rsp_bits_addr; // @[pipe.scala 93:16]
  assign control_io_wid = io_icache_rsp_bits_warpid; // @[pipe.scala 95:17]
  assign operand_collector_clock = clock;
  assign operand_collector_io_control_inst = ibuffer2issue_io_out_bits_inst; // @[pipe.scala 151:31]
  assign operand_collector_io_control_wid = ibuffer2issue_io_out_bits_wid; // @[pipe.scala 151:31]
  assign operand_collector_io_control_branch = ibuffer2issue_io_out_bits_branch; // @[pipe.scala 151:31]
  assign operand_collector_io_control_sel_alu2 = ibuffer2issue_io_out_bits_sel_alu2; // @[pipe.scala 151:31]
  assign operand_collector_io_control_sel_alu1 = ibuffer2issue_io_out_bits_sel_alu1; // @[pipe.scala 151:31]
  assign operand_collector_io_control_isvec = ibuffer2issue_io_out_bits_isvec; // @[pipe.scala 151:31]
  assign operand_collector_io_control_sel_alu3 = ibuffer2issue_io_out_bits_sel_alu3; // @[pipe.scala 151:31]
  assign operand_collector_io_control_mask = ibuffer2issue_io_out_bits_mask; // @[pipe.scala 151:31]
  assign operand_collector_io_control_sel_imm = ibuffer2issue_io_out_bits_sel_imm; // @[pipe.scala 151:31]
  assign operand_collector_io_control_reg_idx1 = ibuffer2issue_io_out_bits_reg_idx1; // @[pipe.scala 151:31]
  assign operand_collector_io_control_reg_idx2 = ibuffer2issue_io_out_bits_reg_idx2; // @[pipe.scala 151:31]
  assign operand_collector_io_control_reg_idx3 = ibuffer2issue_io_out_bits_reg_idx3; // @[pipe.scala 151:31]
  assign operand_collector_io_control_pc = ibuffer2issue_io_out_bits_pc; // @[pipe.scala 151:31]
  assign operand_collector_io_writeScalarCtrl_valid = wb_io_out_x_valid; // @[pipe.scala 153:39]
  assign operand_collector_io_writeScalarCtrl_bits_wb_wxd_rd = wb_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 153:39]
  assign operand_collector_io_writeScalarCtrl_bits_wxd = wb_io_out_x_bits_wxd; // @[pipe.scala 153:39]
  assign operand_collector_io_writeScalarCtrl_bits_reg_idxw = wb_io_out_x_bits_reg_idxw; // @[pipe.scala 153:39]
  assign operand_collector_io_writeScalarCtrl_bits_warp_id = wb_io_out_x_bits_warp_id; // @[pipe.scala 153:39]
  assign operand_collector_io_writeVecCtrl_valid = wb_io_out_v_valid; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_0 = wb_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_1 = wb_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_2 = wb_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_3 = wb_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_4 = wb_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_5 = wb_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_6 = wb_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wb_wfd_rd_7 = wb_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_0 = wb_io_out_v_bits_wfd_mask_0; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_1 = wb_io_out_v_bits_wfd_mask_1; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_2 = wb_io_out_v_bits_wfd_mask_2; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_3 = wb_io_out_v_bits_wfd_mask_3; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_4 = wb_io_out_v_bits_wfd_mask_4; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_5 = wb_io_out_v_bits_wfd_mask_5; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_6 = wb_io_out_v_bits_wfd_mask_6; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd_mask_7 = wb_io_out_v_bits_wfd_mask_7; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_wfd = wb_io_out_v_bits_wfd; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_reg_idxw = wb_io_out_v_bits_reg_idxw; // @[pipe.scala 152:36]
  assign operand_collector_io_writeVecCtrl_bits_warp_id = wb_io_out_v_bits_warp_id; // @[pipe.scala 152:36]
  assign issue_io_in_valid = exe_data_io_deq_valid; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_0 = exe_data_io_deq_bits_in1_0; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_1 = exe_data_io_deq_bits_in1_1; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_2 = exe_data_io_deq_bits_in1_2; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_3 = exe_data_io_deq_bits_in1_3; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_4 = exe_data_io_deq_bits_in1_4; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_5 = exe_data_io_deq_bits_in1_5; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_6 = exe_data_io_deq_bits_in1_6; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in1_7 = exe_data_io_deq_bits_in1_7; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_0 = exe_data_io_deq_bits_in2_0; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_1 = exe_data_io_deq_bits_in2_1; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_2 = exe_data_io_deq_bits_in2_2; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_3 = exe_data_io_deq_bits_in2_3; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_4 = exe_data_io_deq_bits_in2_4; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_5 = exe_data_io_deq_bits_in2_5; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_6 = exe_data_io_deq_bits_in2_6; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in2_7 = exe_data_io_deq_bits_in2_7; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_0 = exe_data_io_deq_bits_in3_0; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_1 = exe_data_io_deq_bits_in3_1; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_2 = exe_data_io_deq_bits_in3_2; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_3 = exe_data_io_deq_bits_in3_3; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_4 = exe_data_io_deq_bits_in3_4; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_5 = exe_data_io_deq_bits_in3_5; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_6 = exe_data_io_deq_bits_in3_6; // @[pipe.scala 214:14]
  assign issue_io_in_bits_in3_7 = exe_data_io_deq_bits_in3_7; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_0 = exe_data_io_deq_bits_mask_0; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_1 = exe_data_io_deq_bits_mask_1; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_2 = exe_data_io_deq_bits_mask_2; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_3 = exe_data_io_deq_bits_mask_3; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_4 = exe_data_io_deq_bits_mask_4; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_5 = exe_data_io_deq_bits_mask_5; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_6 = exe_data_io_deq_bits_mask_6; // @[pipe.scala 214:14]
  assign issue_io_in_bits_mask_7 = exe_data_io_deq_bits_mask_7; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_inst = exe_data_io_deq_bits_ctrl_inst; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_wid = exe_data_io_deq_bits_ctrl_wid; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_fp = exe_data_io_deq_bits_ctrl_fp; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_branch = exe_data_io_deq_bits_ctrl_branch; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_simt_stack = exe_data_io_deq_bits_ctrl_simt_stack; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_simt_stack_op = exe_data_io_deq_bits_ctrl_simt_stack_op; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_barrier = exe_data_io_deq_bits_ctrl_barrier; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_csr = exe_data_io_deq_bits_ctrl_csr; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_reverse = exe_data_io_deq_bits_ctrl_reverse; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_isvec = exe_data_io_deq_bits_ctrl_isvec; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_mem_unsigned = exe_data_io_deq_bits_ctrl_mem_unsigned; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_alu_fn = exe_data_io_deq_bits_ctrl_alu_fn; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_mem = exe_data_io_deq_bits_ctrl_mem; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_mem_cmd = exe_data_io_deq_bits_ctrl_mem_cmd; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_mop = exe_data_io_deq_bits_ctrl_mop; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_reg_idxw = exe_data_io_deq_bits_ctrl_reg_idxw; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_wfd = exe_data_io_deq_bits_ctrl_wfd; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_fence = exe_data_io_deq_bits_ctrl_fence; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_sfu = exe_data_io_deq_bits_ctrl_sfu; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_readmask = exe_data_io_deq_bits_ctrl_readmask; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_writemask = exe_data_io_deq_bits_ctrl_writemask; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_wxd = exe_data_io_deq_bits_ctrl_wxd; // @[pipe.scala 214:14]
  assign issue_io_in_bits_ctrl_pc = exe_data_io_deq_bits_ctrl_pc; // @[pipe.scala 214:14]
  assign issue_io_out_sALU_ready = alu_io_in_ready; // @[pipe.scala 218:20]
  assign issue_io_out_vALU_ready = valu_io_in_ready; // @[pipe.scala 216:20]
  assign issue_io_out_vFPU_ready = fpu_io_in_ready; // @[pipe.scala 228:20]
  assign issue_io_out_LSU_ready = lsu_io_lsu_req_ready; // @[pipe.scala 217:19]
  assign issue_io_out_SFU_ready = sfu_io_in_ready; // @[pipe.scala 221:19]
  assign issue_io_out_SIMT_ready = simt_stack_io_branch_ctl_ready; // @[pipe.scala 220:20]
  assign issue_io_out_warpscheduler_ready = warp_sche_io_warp_control_ready; // @[pipe.scala 74:28]
  assign issue_io_out_CSR_ready = csrfile_io_in_ready; // @[pipe.scala 219:19]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = issue_io_out_sALU_valid; // @[pipe.scala 218:20]
  assign alu_io_in_bits_in1 = issue_io_out_sALU_bits_in1; // @[pipe.scala 218:20]
  assign alu_io_in_bits_in2 = issue_io_out_sALU_bits_in2; // @[pipe.scala 218:20]
  assign alu_io_in_bits_in3 = issue_io_out_sALU_bits_in3; // @[pipe.scala 218:20]
  assign alu_io_in_bits_ctrl_wid = issue_io_out_sALU_bits_ctrl_wid; // @[pipe.scala 218:20]
  assign alu_io_in_bits_ctrl_branch = issue_io_out_sALU_bits_ctrl_branch; // @[pipe.scala 218:20]
  assign alu_io_in_bits_ctrl_alu_fn = issue_io_out_sALU_bits_ctrl_alu_fn; // @[pipe.scala 218:20]
  assign alu_io_in_bits_ctrl_reg_idxw = issue_io_out_sALU_bits_ctrl_reg_idxw; // @[pipe.scala 218:20]
  assign alu_io_in_bits_ctrl_wxd = issue_io_out_sALU_bits_ctrl_wxd; // @[pipe.scala 218:20]
  assign alu_io_out2br_ready = branch_back_io_in0_ready; // @[pipe.scala 226:16]
  assign valu_clock = clock;
  assign valu_reset = reset;
  assign valu_io_in_valid = issue_io_out_vALU_valid; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_0 = issue_io_out_vALU_bits_in1_0; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_1 = issue_io_out_vALU_bits_in1_1; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_2 = issue_io_out_vALU_bits_in1_2; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_3 = issue_io_out_vALU_bits_in1_3; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_4 = issue_io_out_vALU_bits_in1_4; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_5 = issue_io_out_vALU_bits_in1_5; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_6 = issue_io_out_vALU_bits_in1_6; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in1_7 = issue_io_out_vALU_bits_in1_7; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_0 = issue_io_out_vALU_bits_in2_0; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_1 = issue_io_out_vALU_bits_in2_1; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_2 = issue_io_out_vALU_bits_in2_2; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_3 = issue_io_out_vALU_bits_in2_3; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_4 = issue_io_out_vALU_bits_in2_4; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_5 = issue_io_out_vALU_bits_in2_5; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_6 = issue_io_out_vALU_bits_in2_6; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in2_7 = issue_io_out_vALU_bits_in2_7; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_0 = issue_io_out_vALU_bits_in3_0; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_1 = issue_io_out_vALU_bits_in3_1; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_2 = issue_io_out_vALU_bits_in3_2; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_3 = issue_io_out_vALU_bits_in3_3; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_4 = issue_io_out_vALU_bits_in3_4; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_5 = issue_io_out_vALU_bits_in3_5; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_6 = issue_io_out_vALU_bits_in3_6; // @[pipe.scala 216:20]
  assign valu_io_in_bits_in3_7 = issue_io_out_vALU_bits_in3_7; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_0 = issue_io_out_vALU_bits_mask_0; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_1 = issue_io_out_vALU_bits_mask_1; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_2 = issue_io_out_vALU_bits_mask_2; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_3 = issue_io_out_vALU_bits_mask_3; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_4 = issue_io_out_vALU_bits_mask_4; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_5 = issue_io_out_vALU_bits_mask_5; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_6 = issue_io_out_vALU_bits_mask_6; // @[pipe.scala 216:20]
  assign valu_io_in_bits_mask_7 = issue_io_out_vALU_bits_mask_7; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_wid = issue_io_out_vALU_bits_ctrl_wid; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_simt_stack = issue_io_out_vALU_bits_ctrl_simt_stack; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_reverse = issue_io_out_vALU_bits_ctrl_reverse; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_alu_fn = issue_io_out_vALU_bits_ctrl_alu_fn; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_reg_idxw = issue_io_out_vALU_bits_ctrl_reg_idxw; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_wfd = issue_io_out_vALU_bits_ctrl_wfd; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_readmask = issue_io_out_vALU_bits_ctrl_readmask; // @[pipe.scala 216:20]
  assign valu_io_in_bits_ctrl_writemask = issue_io_out_vALU_bits_ctrl_writemask; // @[pipe.scala 216:20]
  assign valu_io_out2simt_stack_ready = simt_stack_io_if_mask_ready; // @[pipe.scala 223:24]
  assign fpu_clock = clock;
  assign fpu_reset = reset;
  assign fpu_io_in_valid = issue_io_out_vFPU_valid; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_0 = issue_io_out_vFPU_bits_in1_0; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_1 = issue_io_out_vFPU_bits_in1_1; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_2 = issue_io_out_vFPU_bits_in1_2; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_3 = issue_io_out_vFPU_bits_in1_3; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_4 = issue_io_out_vFPU_bits_in1_4; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_5 = issue_io_out_vFPU_bits_in1_5; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_6 = issue_io_out_vFPU_bits_in1_6; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in1_7 = issue_io_out_vFPU_bits_in1_7; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_0 = issue_io_out_vFPU_bits_in2_0; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_1 = issue_io_out_vFPU_bits_in2_1; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_2 = issue_io_out_vFPU_bits_in2_2; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_3 = issue_io_out_vFPU_bits_in2_3; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_4 = issue_io_out_vFPU_bits_in2_4; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_5 = issue_io_out_vFPU_bits_in2_5; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_6 = issue_io_out_vFPU_bits_in2_6; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in2_7 = issue_io_out_vFPU_bits_in2_7; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_0 = issue_io_out_vFPU_bits_in3_0; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_1 = issue_io_out_vFPU_bits_in3_1; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_2 = issue_io_out_vFPU_bits_in3_2; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_3 = issue_io_out_vFPU_bits_in3_3; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_4 = issue_io_out_vFPU_bits_in3_4; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_5 = issue_io_out_vFPU_bits_in3_5; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_6 = issue_io_out_vFPU_bits_in3_6; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_in3_7 = issue_io_out_vFPU_bits_in3_7; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_0 = issue_io_out_vFPU_bits_mask_0; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_1 = issue_io_out_vFPU_bits_mask_1; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_2 = issue_io_out_vFPU_bits_mask_2; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_3 = issue_io_out_vFPU_bits_mask_3; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_4 = issue_io_out_vFPU_bits_mask_4; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_5 = issue_io_out_vFPU_bits_mask_5; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_6 = issue_io_out_vFPU_bits_mask_6; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_mask_7 = issue_io_out_vFPU_bits_mask_7; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_ctrl_wid = issue_io_out_vFPU_bits_ctrl_wid; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_ctrl_reverse = issue_io_out_vFPU_bits_ctrl_reverse; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_ctrl_alu_fn = issue_io_out_vFPU_bits_ctrl_alu_fn; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_ctrl_reg_idxw = issue_io_out_vFPU_bits_ctrl_reg_idxw; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_ctrl_wfd = issue_io_out_vFPU_bits_ctrl_wfd; // @[pipe.scala 228:20]
  assign fpu_io_in_bits_ctrl_wxd = issue_io_out_vFPU_bits_ctrl_wxd; // @[pipe.scala 228:20]
  assign fpu_io_rm = csrfile_io_frm; // @[pipe.scala 229:12]
  assign fpu_io_out_x_ready = wb_io_in_x_1_ready; // @[pipe.scala 240:16]
  assign fpu_io_out_v_ready = wb_io_in_v_1_ready; // @[pipe.scala 245:16]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_lsu_req_valid = issue_io_out_LSU_valid; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_0 = issue_io_out_LSU_bits_in1_0; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_1 = issue_io_out_LSU_bits_in1_1; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_2 = issue_io_out_LSU_bits_in1_2; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_3 = issue_io_out_LSU_bits_in1_3; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_4 = issue_io_out_LSU_bits_in1_4; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_5 = issue_io_out_LSU_bits_in1_5; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_6 = issue_io_out_LSU_bits_in1_6; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in1_7 = issue_io_out_LSU_bits_in1_7; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_0 = issue_io_out_LSU_bits_in2_0; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_1 = issue_io_out_LSU_bits_in2_1; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_2 = issue_io_out_LSU_bits_in2_2; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_3 = issue_io_out_LSU_bits_in2_3; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_4 = issue_io_out_LSU_bits_in2_4; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_5 = issue_io_out_LSU_bits_in2_5; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_6 = issue_io_out_LSU_bits_in2_6; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in2_7 = issue_io_out_LSU_bits_in2_7; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_0 = issue_io_out_LSU_bits_in3_0; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_1 = issue_io_out_LSU_bits_in3_1; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_2 = issue_io_out_LSU_bits_in3_2; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_3 = issue_io_out_LSU_bits_in3_3; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_4 = issue_io_out_LSU_bits_in3_4; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_5 = issue_io_out_LSU_bits_in3_5; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_6 = issue_io_out_LSU_bits_in3_6; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_in3_7 = issue_io_out_LSU_bits_in3_7; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_0 = issue_io_out_LSU_bits_mask_0; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_1 = issue_io_out_LSU_bits_mask_1; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_2 = issue_io_out_LSU_bits_mask_2; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_3 = issue_io_out_LSU_bits_mask_3; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_4 = issue_io_out_LSU_bits_mask_4; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_5 = issue_io_out_LSU_bits_mask_5; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_6 = issue_io_out_LSU_bits_mask_6; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_mask_7 = issue_io_out_LSU_bits_mask_7; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_inst = issue_io_out_LSU_bits_ctrl_inst; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_wid = issue_io_out_LSU_bits_ctrl_wid; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_fp = issue_io_out_LSU_bits_ctrl_fp; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_branch = issue_io_out_LSU_bits_ctrl_branch; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_simt_stack = issue_io_out_LSU_bits_ctrl_simt_stack; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_simt_stack_op = issue_io_out_LSU_bits_ctrl_simt_stack_op; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_barrier = issue_io_out_LSU_bits_ctrl_barrier; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_csr = issue_io_out_LSU_bits_ctrl_csr; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_reverse = issue_io_out_LSU_bits_ctrl_reverse; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_isvec = issue_io_out_LSU_bits_ctrl_isvec; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_mem_unsigned = issue_io_out_LSU_bits_ctrl_mem_unsigned; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_alu_fn = issue_io_out_LSU_bits_ctrl_alu_fn; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_mem = issue_io_out_LSU_bits_ctrl_mem; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_mem_cmd = issue_io_out_LSU_bits_ctrl_mem_cmd; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_mop = issue_io_out_LSU_bits_ctrl_mop; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_reg_idxw = issue_io_out_LSU_bits_ctrl_reg_idxw; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_wfd = issue_io_out_LSU_bits_ctrl_wfd; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_fence = issue_io_out_LSU_bits_ctrl_fence; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_sfu = issue_io_out_LSU_bits_ctrl_sfu; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_readmask = issue_io_out_LSU_bits_ctrl_readmask; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_writemask = issue_io_out_LSU_bits_ctrl_writemask; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_wxd = issue_io_out_LSU_bits_ctrl_wxd; // @[pipe.scala 217:19]
  assign lsu_io_lsu_req_bits_ctrl_pc = issue_io_out_LSU_bits_ctrl_pc; // @[pipe.scala 217:19]
  assign lsu_io_dcache_rsp_valid = io_dcache_rsp_valid; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_instrId = io_dcache_rsp_bits_instrId; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_0 = io_dcache_rsp_bits_data_0; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_1 = io_dcache_rsp_bits_data_1; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_2 = io_dcache_rsp_bits_data_2; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_3 = io_dcache_rsp_bits_data_3; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_4 = io_dcache_rsp_bits_data_4; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_5 = io_dcache_rsp_bits_data_5; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_6 = io_dcache_rsp_bits_data_6; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_data_7 = io_dcache_rsp_bits_data_7; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_0 = io_dcache_rsp_bits_activeMask_0; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_1 = io_dcache_rsp_bits_activeMask_1; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_2 = io_dcache_rsp_bits_activeMask_2; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_3 = io_dcache_rsp_bits_activeMask_3; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_4 = io_dcache_rsp_bits_activeMask_4; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_5 = io_dcache_rsp_bits_activeMask_5; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_6 = io_dcache_rsp_bits_activeMask_6; // @[pipe.scala 233:20]
  assign lsu_io_dcache_rsp_bits_activeMask_7 = io_dcache_rsp_bits_activeMask_7; // @[pipe.scala 233:20]
  assign lsu_io_lsu_rsp_ready = lsu2wb_io_lsu_rsp_ready; // @[pipe.scala 235:17]
  assign lsu_io_dcache_req_ready = io_dcache_req_ready; // @[pipe.scala 234:20]
  assign lsu_io_shared_req_ready = io_shared_req_ready; // @[pipe.scala 237:20]
  assign lsu_io_shared_rsp_valid = io_shared_rsp_valid; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_instrId = io_shared_rsp_bits_instrId; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_0 = io_shared_rsp_bits_data_0; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_1 = io_shared_rsp_bits_data_1; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_2 = io_shared_rsp_bits_data_2; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_3 = io_shared_rsp_bits_data_3; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_4 = io_shared_rsp_bits_data_4; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_5 = io_shared_rsp_bits_data_5; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_6 = io_shared_rsp_bits_data_6; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_data_7 = io_shared_rsp_bits_data_7; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_0 = io_shared_rsp_bits_activeMask_0; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_1 = io_shared_rsp_bits_activeMask_1; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_2 = io_shared_rsp_bits_activeMask_2; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_3 = io_shared_rsp_bits_activeMask_3; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_4 = io_shared_rsp_bits_activeMask_4; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_5 = io_shared_rsp_bits_activeMask_5; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_6 = io_shared_rsp_bits_activeMask_6; // @[pipe.scala 236:20]
  assign lsu_io_shared_rsp_bits_activeMask_7 = io_shared_rsp_bits_activeMask_7; // @[pipe.scala 236:20]
  assign sfu_clock = clock;
  assign sfu_reset = reset;
  assign sfu_io_in_valid = issue_io_out_SFU_valid; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_0 = issue_io_out_SFU_bits_in1_0; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_1 = issue_io_out_SFU_bits_in1_1; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_2 = issue_io_out_SFU_bits_in1_2; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_3 = issue_io_out_SFU_bits_in1_3; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_4 = issue_io_out_SFU_bits_in1_4; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_5 = issue_io_out_SFU_bits_in1_5; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_6 = issue_io_out_SFU_bits_in1_6; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in1_7 = issue_io_out_SFU_bits_in1_7; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_0 = issue_io_out_SFU_bits_in2_0; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_1 = issue_io_out_SFU_bits_in2_1; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_2 = issue_io_out_SFU_bits_in2_2; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_3 = issue_io_out_SFU_bits_in2_3; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_4 = issue_io_out_SFU_bits_in2_4; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_5 = issue_io_out_SFU_bits_in2_5; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_6 = issue_io_out_SFU_bits_in2_6; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_in2_7 = issue_io_out_SFU_bits_in2_7; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_0 = issue_io_out_SFU_bits_mask_0; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_1 = issue_io_out_SFU_bits_mask_1; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_2 = issue_io_out_SFU_bits_mask_2; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_3 = issue_io_out_SFU_bits_mask_3; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_4 = issue_io_out_SFU_bits_mask_4; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_5 = issue_io_out_SFU_bits_mask_5; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_6 = issue_io_out_SFU_bits_mask_6; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_mask_7 = issue_io_out_SFU_bits_mask_7; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_wid = issue_io_out_SFU_bits_ctrl_wid; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_fp = issue_io_out_SFU_bits_ctrl_fp; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_reverse = issue_io_out_SFU_bits_ctrl_reverse; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_isvec = issue_io_out_SFU_bits_ctrl_isvec; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_alu_fn = issue_io_out_SFU_bits_ctrl_alu_fn; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_reg_idxw = issue_io_out_SFU_bits_ctrl_reg_idxw; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_wfd = issue_io_out_SFU_bits_ctrl_wfd; // @[pipe.scala 221:19]
  assign sfu_io_in_bits_ctrl_wxd = issue_io_out_SFU_bits_ctrl_wxd; // @[pipe.scala 221:19]
  assign sfu_io_rm = csrfile_io_frm; // @[pipe.scala 230:12]
  assign sfu_io_out_x_ready = wb_io_in_x_4_ready; // @[pipe.scala 243:16]
  assign sfu_io_out_v_ready = wb_io_in_v_3_ready; // @[pipe.scala 247:16]
  assign lsu2wb_io_lsu_rsp_valid = lsu_io_lsu_rsp_valid; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_warp_id = lsu_io_lsu_rsp_bits_tag_warp_id; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_wfd = lsu_io_lsu_rsp_bits_tag_wfd; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_wxd = lsu_io_lsu_rsp_bits_tag_wxd; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_reg_idxw = lsu_io_lsu_rsp_bits_tag_reg_idxw; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_0 = lsu_io_lsu_rsp_bits_tag_mask_0; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_1 = lsu_io_lsu_rsp_bits_tag_mask_1; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_2 = lsu_io_lsu_rsp_bits_tag_mask_2; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_3 = lsu_io_lsu_rsp_bits_tag_mask_3; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_4 = lsu_io_lsu_rsp_bits_tag_mask_4; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_5 = lsu_io_lsu_rsp_bits_tag_mask_5; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_6 = lsu_io_lsu_rsp_bits_tag_mask_6; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_mask_7 = lsu_io_lsu_rsp_bits_tag_mask_7; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_tag_isWrite = lsu_io_lsu_rsp_bits_tag_isWrite; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_0 = lsu_io_lsu_rsp_bits_data_0; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_1 = lsu_io_lsu_rsp_bits_data_1; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_2 = lsu_io_lsu_rsp_bits_data_2; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_3 = lsu_io_lsu_rsp_bits_data_3; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_4 = lsu_io_lsu_rsp_bits_data_4; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_5 = lsu_io_lsu_rsp_bits_data_5; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_6 = lsu_io_lsu_rsp_bits_data_6; // @[pipe.scala 235:17]
  assign lsu2wb_io_lsu_rsp_bits_data_7 = lsu_io_lsu_rsp_bits_data_7; // @[pipe.scala 235:17]
  assign lsu2wb_io_out_x_ready = wb_io_in_x_2_ready; // @[pipe.scala 241:16]
  assign lsu2wb_io_out_v_ready = wb_io_in_v_2_ready; // @[pipe.scala 246:16]
  assign wb_io_out_v_ready = 1'h1; // @[pipe.scala 152:36]
  assign wb_io_out_x_ready = 1'h1; // @[pipe.scala 153:39]
  assign wb_io_in_x_0_valid = alu_io_out_valid; // @[pipe.scala 239:16]
  assign wb_io_in_x_0_bits_wb_wxd_rd = alu_io_out_bits_wb_wxd_rd; // @[pipe.scala 239:16]
  assign wb_io_in_x_0_bits_wxd = alu_io_out_bits_wxd; // @[pipe.scala 239:16]
  assign wb_io_in_x_0_bits_reg_idxw = alu_io_out_bits_reg_idxw; // @[pipe.scala 239:16]
  assign wb_io_in_x_0_bits_warp_id = alu_io_out_bits_warp_id; // @[pipe.scala 239:16]
  assign wb_io_in_x_1_valid = fpu_io_out_x_valid; // @[pipe.scala 240:16]
  assign wb_io_in_x_1_bits_wb_wxd_rd = fpu_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 240:16]
  assign wb_io_in_x_1_bits_wxd = fpu_io_out_x_bits_wxd; // @[pipe.scala 240:16]
  assign wb_io_in_x_1_bits_reg_idxw = fpu_io_out_x_bits_reg_idxw; // @[pipe.scala 240:16]
  assign wb_io_in_x_1_bits_warp_id = fpu_io_out_x_bits_warp_id; // @[pipe.scala 240:16]
  assign wb_io_in_x_2_valid = lsu2wb_io_out_x_valid; // @[pipe.scala 241:16]
  assign wb_io_in_x_2_bits_wb_wxd_rd = lsu2wb_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 241:16]
  assign wb_io_in_x_2_bits_wxd = lsu2wb_io_out_x_bits_wxd; // @[pipe.scala 241:16]
  assign wb_io_in_x_2_bits_reg_idxw = lsu2wb_io_out_x_bits_reg_idxw; // @[pipe.scala 241:16]
  assign wb_io_in_x_2_bits_warp_id = lsu2wb_io_out_x_bits_warp_id; // @[pipe.scala 241:16]
  assign wb_io_in_x_3_valid = csrfile_io_out_valid; // @[pipe.scala 242:16]
  assign wb_io_in_x_3_bits_wb_wxd_rd = csrfile_io_out_bits_wb_wxd_rd; // @[pipe.scala 242:16]
  assign wb_io_in_x_3_bits_wxd = csrfile_io_out_bits_wxd; // @[pipe.scala 242:16]
  assign wb_io_in_x_3_bits_reg_idxw = csrfile_io_out_bits_reg_idxw; // @[pipe.scala 242:16]
  assign wb_io_in_x_3_bits_warp_id = csrfile_io_out_bits_warp_id; // @[pipe.scala 242:16]
  assign wb_io_in_x_4_valid = sfu_io_out_x_valid; // @[pipe.scala 243:16]
  assign wb_io_in_x_4_bits_wb_wxd_rd = sfu_io_out_x_bits_wb_wxd_rd; // @[pipe.scala 243:16]
  assign wb_io_in_x_4_bits_wxd = sfu_io_out_x_bits_wxd; // @[pipe.scala 243:16]
  assign wb_io_in_x_4_bits_reg_idxw = sfu_io_out_x_bits_reg_idxw; // @[pipe.scala 243:16]
  assign wb_io_in_x_4_bits_warp_id = sfu_io_out_x_bits_warp_id; // @[pipe.scala 243:16]
  assign wb_io_in_v_0_valid = valu_io_out_valid; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_0 = valu_io_out_bits_wb_wfd_rd_0; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_1 = valu_io_out_bits_wb_wfd_rd_1; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_2 = valu_io_out_bits_wb_wfd_rd_2; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_3 = valu_io_out_bits_wb_wfd_rd_3; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_4 = valu_io_out_bits_wb_wfd_rd_4; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_5 = valu_io_out_bits_wb_wfd_rd_5; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_6 = valu_io_out_bits_wb_wfd_rd_6; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wb_wfd_rd_7 = valu_io_out_bits_wb_wfd_rd_7; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_0 = valu_io_out_bits_wfd_mask_0; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_1 = valu_io_out_bits_wfd_mask_1; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_2 = valu_io_out_bits_wfd_mask_2; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_3 = valu_io_out_bits_wfd_mask_3; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_4 = valu_io_out_bits_wfd_mask_4; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_5 = valu_io_out_bits_wfd_mask_5; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_6 = valu_io_out_bits_wfd_mask_6; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd_mask_7 = valu_io_out_bits_wfd_mask_7; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_wfd = valu_io_out_bits_wfd; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_reg_idxw = valu_io_out_bits_reg_idxw; // @[pipe.scala 244:16]
  assign wb_io_in_v_0_bits_warp_id = valu_io_out_bits_warp_id; // @[pipe.scala 244:16]
  assign wb_io_in_v_1_valid = fpu_io_out_v_valid; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_0 = fpu_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_1 = fpu_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_2 = fpu_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_3 = fpu_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_4 = fpu_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_5 = fpu_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_6 = fpu_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wb_wfd_rd_7 = fpu_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_0 = fpu_io_out_v_bits_wfd_mask_0; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_1 = fpu_io_out_v_bits_wfd_mask_1; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_2 = fpu_io_out_v_bits_wfd_mask_2; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_3 = fpu_io_out_v_bits_wfd_mask_3; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_4 = fpu_io_out_v_bits_wfd_mask_4; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_5 = fpu_io_out_v_bits_wfd_mask_5; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_6 = fpu_io_out_v_bits_wfd_mask_6; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd_mask_7 = fpu_io_out_v_bits_wfd_mask_7; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_wfd = fpu_io_out_v_bits_wfd; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_reg_idxw = fpu_io_out_v_bits_reg_idxw; // @[pipe.scala 245:16]
  assign wb_io_in_v_1_bits_warp_id = fpu_io_out_v_bits_warp_id; // @[pipe.scala 245:16]
  assign wb_io_in_v_2_valid = lsu2wb_io_out_v_valid; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_0 = lsu2wb_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_1 = lsu2wb_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_2 = lsu2wb_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_3 = lsu2wb_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_4 = lsu2wb_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_5 = lsu2wb_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_6 = lsu2wb_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wb_wfd_rd_7 = lsu2wb_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_0 = lsu2wb_io_out_v_bits_wfd_mask_0; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_1 = lsu2wb_io_out_v_bits_wfd_mask_1; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_2 = lsu2wb_io_out_v_bits_wfd_mask_2; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_3 = lsu2wb_io_out_v_bits_wfd_mask_3; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_4 = lsu2wb_io_out_v_bits_wfd_mask_4; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_5 = lsu2wb_io_out_v_bits_wfd_mask_5; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_6 = lsu2wb_io_out_v_bits_wfd_mask_6; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd_mask_7 = lsu2wb_io_out_v_bits_wfd_mask_7; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_wfd = lsu2wb_io_out_v_bits_wfd; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_reg_idxw = lsu2wb_io_out_v_bits_reg_idxw; // @[pipe.scala 246:16]
  assign wb_io_in_v_2_bits_warp_id = lsu2wb_io_out_v_bits_warp_id; // @[pipe.scala 246:16]
  assign wb_io_in_v_3_valid = sfu_io_out_v_valid; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_0 = sfu_io_out_v_bits_wb_wfd_rd_0; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_1 = sfu_io_out_v_bits_wb_wfd_rd_1; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_2 = sfu_io_out_v_bits_wb_wfd_rd_2; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_3 = sfu_io_out_v_bits_wb_wfd_rd_3; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_4 = sfu_io_out_v_bits_wb_wfd_rd_4; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_5 = sfu_io_out_v_bits_wb_wfd_rd_5; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_6 = sfu_io_out_v_bits_wb_wfd_rd_6; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wb_wfd_rd_7 = sfu_io_out_v_bits_wb_wfd_rd_7; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_0 = sfu_io_out_v_bits_wfd_mask_0; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_1 = sfu_io_out_v_bits_wfd_mask_1; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_2 = sfu_io_out_v_bits_wfd_mask_2; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_3 = sfu_io_out_v_bits_wfd_mask_3; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_4 = sfu_io_out_v_bits_wfd_mask_4; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_5 = sfu_io_out_v_bits_wfd_mask_5; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_6 = sfu_io_out_v_bits_wfd_mask_6; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd_mask_7 = sfu_io_out_v_bits_wfd_mask_7; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_wfd = sfu_io_out_v_bits_wfd; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_reg_idxw = sfu_io_out_v_bits_reg_idxw; // @[pipe.scala 247:16]
  assign wb_io_in_v_3_bits_warp_id = sfu_io_out_v_bits_warp_id; // @[pipe.scala 247:16]
  assign Scoreboard_clock = clock;
  assign Scoreboard_reset = reset;
  assign Scoreboard_io_ibuffer_if_ctrl_sel_alu2 = ibuffer_io_out_0_bits_sel_alu2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_sel_alu1 = ibuffer_io_out_0_bits_sel_alu1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_isvec = ibuffer_io_out_0_bits_isvec; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_sel_alu3 = ibuffer_io_out_0_bits_sel_alu3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_mask = ibuffer_io_out_0_bits_mask; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_mem = ibuffer_io_out_0_bits_mem; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_reg_idx1 = ibuffer_io_out_0_bits_reg_idx1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_reg_idx2 = ibuffer_io_out_0_bits_reg_idx2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_ibuffer_if_ctrl_reg_idx3 = ibuffer_io_out_0_bits_reg_idx3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_io_if_ctrl_branch = exe_data_io_enq_bits_ctrl_branch; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_io_if_ctrl_barrier = exe_data_io_enq_bits_ctrl_barrier; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_io_if_ctrl_reg_idxw = exe_data_io_enq_bits_ctrl_reg_idxw; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_io_if_ctrl_wfd = exe_data_io_enq_bits_ctrl_wfd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_io_if_ctrl_fence = exe_data_io_enq_bits_ctrl_fence; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_io_if_ctrl_wxd = exe_data_io_enq_bits_ctrl_wxd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_io_wb_v_ctrl_wfd = wb_io_out_v_bits_wfd; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_io_wb_v_ctrl_reg_idxw = wb_io_out_v_bits_reg_idxw; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_io_wb_x_ctrl_wxd = wb_io_out_x_bits_wxd; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_io_wb_x_ctrl_reg_idxw = wb_io_out_x_bits_reg_idxw; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_io_if_fire = 2'h0 == exe_data_io_enq_bits_ctrl_wid & _warp_sche_io_issued_warp_valid_T; // @[pipe.scala 139:22 147:{48,48}]
  assign Scoreboard_io_br_ctrl = _T_4 & warp_sche_io_branch_bits_wid == 2'h0 | _GEN_1; // @[pipe.scala 143:{81,99}]
  assign Scoreboard_io_fence_end = lsu_io_fence_end[0]; // @[pipe.scala 138:42]
  assign Scoreboard_io_wb_v_fire = 2'h0 == wb_io_out_v_bits_warp_id & _scoreb_wb_v_fire_T; // @[pipe.scala 140:24 149:{45,45}]
  assign Scoreboard_io_wb_x_fire = 2'h0 == wb_io_out_x_bits_warp_id & _scoreb_wb_x_fire_T; // @[pipe.scala 141:24 148:{45,45}]
  assign Scoreboard_1_clock = clock;
  assign Scoreboard_1_reset = reset;
  assign Scoreboard_1_io_ibuffer_if_ctrl_sel_alu2 = ibuffer_io_out_1_bits_sel_alu2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_sel_alu1 = ibuffer_io_out_1_bits_sel_alu1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_isvec = ibuffer_io_out_1_bits_isvec; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_sel_alu3 = ibuffer_io_out_1_bits_sel_alu3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_mask = ibuffer_io_out_1_bits_mask; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_mem = ibuffer_io_out_1_bits_mem; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_reg_idx1 = ibuffer_io_out_1_bits_reg_idx1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_reg_idx2 = ibuffer_io_out_1_bits_reg_idx2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_ibuffer_if_ctrl_reg_idx3 = ibuffer_io_out_1_bits_reg_idx3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_1_io_if_ctrl_branch = exe_data_io_enq_bits_ctrl_branch; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_1_io_if_ctrl_barrier = exe_data_io_enq_bits_ctrl_barrier; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_1_io_if_ctrl_reg_idxw = exe_data_io_enq_bits_ctrl_reg_idxw; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_1_io_if_ctrl_wfd = exe_data_io_enq_bits_ctrl_wfd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_1_io_if_ctrl_fence = exe_data_io_enq_bits_ctrl_fence; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_1_io_if_ctrl_wxd = exe_data_io_enq_bits_ctrl_wxd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_1_io_wb_v_ctrl_wfd = wb_io_out_v_bits_wfd; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_1_io_wb_v_ctrl_reg_idxw = wb_io_out_v_bits_reg_idxw; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_1_io_wb_x_ctrl_wxd = wb_io_out_x_bits_wxd; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_1_io_wb_x_ctrl_reg_idxw = wb_io_out_x_bits_reg_idxw; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_1_io_if_fire = 2'h1 == exe_data_io_enq_bits_ctrl_wid & _warp_sche_io_issued_warp_valid_T; // @[pipe.scala 139:22 147:{48,48}]
  assign Scoreboard_1_io_br_ctrl = _T_4 & warp_sche_io_branch_bits_wid == 2'h1 | _GEN_4; // @[pipe.scala 143:{81,99}]
  assign Scoreboard_1_io_fence_end = lsu_io_fence_end[1]; // @[pipe.scala 138:42]
  assign Scoreboard_1_io_wb_v_fire = 2'h1 == wb_io_out_v_bits_warp_id & _scoreb_wb_v_fire_T; // @[pipe.scala 140:24 149:{45,45}]
  assign Scoreboard_1_io_wb_x_fire = 2'h1 == wb_io_out_x_bits_warp_id & _scoreb_wb_x_fire_T; // @[pipe.scala 141:24 148:{45,45}]
  assign Scoreboard_2_clock = clock;
  assign Scoreboard_2_reset = reset;
  assign Scoreboard_2_io_ibuffer_if_ctrl_sel_alu2 = ibuffer_io_out_2_bits_sel_alu2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_sel_alu1 = ibuffer_io_out_2_bits_sel_alu1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_isvec = ibuffer_io_out_2_bits_isvec; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_sel_alu3 = ibuffer_io_out_2_bits_sel_alu3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_mask = ibuffer_io_out_2_bits_mask; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_mem = ibuffer_io_out_2_bits_mem; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_reg_idx1 = ibuffer_io_out_2_bits_reg_idx1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_reg_idx2 = ibuffer_io_out_2_bits_reg_idx2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_ibuffer_if_ctrl_reg_idx3 = ibuffer_io_out_2_bits_reg_idx3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_2_io_if_ctrl_branch = exe_data_io_enq_bits_ctrl_branch; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_2_io_if_ctrl_barrier = exe_data_io_enq_bits_ctrl_barrier; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_2_io_if_ctrl_reg_idxw = exe_data_io_enq_bits_ctrl_reg_idxw; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_2_io_if_ctrl_wfd = exe_data_io_enq_bits_ctrl_wfd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_2_io_if_ctrl_fence = exe_data_io_enq_bits_ctrl_fence; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_2_io_if_ctrl_wxd = exe_data_io_enq_bits_ctrl_wxd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_2_io_wb_v_ctrl_wfd = wb_io_out_v_bits_wfd; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_2_io_wb_v_ctrl_reg_idxw = wb_io_out_v_bits_reg_idxw; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_2_io_wb_x_ctrl_wxd = wb_io_out_x_bits_wxd; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_2_io_wb_x_ctrl_reg_idxw = wb_io_out_x_bits_reg_idxw; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_2_io_if_fire = 2'h2 == exe_data_io_enq_bits_ctrl_wid & _warp_sche_io_issued_warp_valid_T; // @[pipe.scala 139:22 147:{48,48}]
  assign Scoreboard_2_io_br_ctrl = _T_4 & warp_sche_io_branch_bits_wid == 2'h2 | _GEN_7; // @[pipe.scala 143:{81,99}]
  assign Scoreboard_2_io_fence_end = lsu_io_fence_end[2]; // @[pipe.scala 138:42]
  assign Scoreboard_2_io_wb_v_fire = 2'h2 == wb_io_out_v_bits_warp_id & _scoreb_wb_v_fire_T; // @[pipe.scala 140:24 149:{45,45}]
  assign Scoreboard_2_io_wb_x_fire = 2'h2 == wb_io_out_x_bits_warp_id & _scoreb_wb_x_fire_T; // @[pipe.scala 141:24 148:{45,45}]
  assign Scoreboard_3_clock = clock;
  assign Scoreboard_3_reset = reset;
  assign Scoreboard_3_io_ibuffer_if_ctrl_sel_alu2 = ibuffer_io_out_3_bits_sel_alu2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_sel_alu1 = ibuffer_io_out_3_bits_sel_alu1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_isvec = ibuffer_io_out_3_bits_isvec; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_sel_alu3 = ibuffer_io_out_3_bits_sel_alu3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_mask = ibuffer_io_out_3_bits_mask; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_mem = ibuffer_io_out_3_bits_mem; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_reg_idx1 = ibuffer_io_out_3_bits_reg_idx1; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_reg_idx2 = ibuffer_io_out_3_bits_reg_idx2; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_ibuffer_if_ctrl_reg_idx3 = ibuffer_io_out_3_bits_reg_idx3; // @[pipe.scala 52:21 134:30]
  assign Scoreboard_3_io_if_ctrl_branch = exe_data_io_enq_bits_ctrl_branch; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_3_io_if_ctrl_barrier = exe_data_io_enq_bits_ctrl_barrier; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_3_io_if_ctrl_reg_idxw = exe_data_io_enq_bits_ctrl_reg_idxw; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_3_io_if_ctrl_wfd = exe_data_io_enq_bits_ctrl_wfd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_3_io_if_ctrl_fence = exe_data_io_enq_bits_ctrl_fence; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_3_io_if_ctrl_wxd = exe_data_io_enq_bits_ctrl_wxd; // @[pipe.scala 52:21 135:22]
  assign Scoreboard_3_io_wb_v_ctrl_wfd = wb_io_out_v_bits_wfd; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_3_io_wb_v_ctrl_reg_idxw = wb_io_out_v_bits_reg_idxw; // @[pipe.scala 52:21 136:24]
  assign Scoreboard_3_io_wb_x_ctrl_wxd = wb_io_out_x_bits_wxd; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_3_io_wb_x_ctrl_reg_idxw = wb_io_out_x_bits_reg_idxw; // @[pipe.scala 52:21 137:24]
  assign Scoreboard_3_io_if_fire = 2'h3 == exe_data_io_enq_bits_ctrl_wid & _warp_sche_io_issued_warp_valid_T; // @[pipe.scala 139:22 147:{48,48}]
  assign Scoreboard_3_io_br_ctrl = _T_4 & warp_sche_io_branch_bits_wid == 2'h3 | _GEN_10; // @[pipe.scala 143:{81,99}]
  assign Scoreboard_3_io_fence_end = lsu_io_fence_end[3]; // @[pipe.scala 138:42]
  assign Scoreboard_3_io_wb_v_fire = 2'h3 == wb_io_out_v_bits_warp_id & _scoreb_wb_v_fire_T; // @[pipe.scala 140:24 149:{45,45}]
  assign Scoreboard_3_io_wb_x_fire = 2'h3 == wb_io_out_x_bits_warp_id & _scoreb_wb_x_fire_T; // @[pipe.scala 141:24 148:{45,45}]
  assign ibuffer_clock = clock;
  assign ibuffer_reset = reset;
  assign ibuffer_io_in_valid = io_icache_rsp_valid & ~io_icache_rsp_bits_status[0]; // @[pipe.scala 98:43]
  assign ibuffer_io_in_bits_inst = control_io_control_inst; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_wid = control_io_control_wid; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_fp = control_io_control_fp; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_branch = control_io_control_branch; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_simt_stack = control_io_control_simt_stack; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_simt_stack_op = control_io_control_simt_stack_op; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_barrier = control_io_control_barrier; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_csr = control_io_control_csr; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_reverse = control_io_control_reverse; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_sel_alu2 = control_io_control_sel_alu2; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_sel_alu1 = control_io_control_sel_alu1; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_isvec = control_io_control_isvec; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_sel_alu3 = control_io_control_sel_alu3; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_mask = control_io_control_mask; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_sel_imm = control_io_control_sel_imm; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_mem_unsigned = control_io_control_mem_unsigned; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_alu_fn = control_io_control_alu_fn; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_mem = control_io_control_mem; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_mem_cmd = control_io_control_mem_cmd; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_mop = control_io_control_mop; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_reg_idx1 = control_io_control_reg_idx1; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_reg_idx2 = control_io_control_reg_idx2; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_reg_idx3 = control_io_control_reg_idx3; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_reg_idxw = control_io_control_reg_idxw; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_wfd = control_io_control_wfd; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_fence = control_io_control_fence; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_sfu = control_io_control_sfu; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_readmask = control_io_control_readmask; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_writemask = control_io_control_writemask; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_wxd = control_io_control_wxd; // @[pipe.scala 97:21]
  assign ibuffer_io_in_bits_pc = control_io_control_pc; // @[pipe.scala 97:21]
  assign ibuffer_io_flush_valid = warp_sche_io_flush_valid; // @[pipe.scala 99:19]
  assign ibuffer_io_flush_bits = warp_sche_io_flush_bits; // @[pipe.scala 99:19]
  assign ibuffer_io_out_0_ready = ibuffer2issue_io_in_0_ready & warp_sche_io_warp_ready[0]; // @[pipe.scala 121:59]
  assign ibuffer_io_out_1_ready = ibuffer2issue_io_in_1_ready & warp_sche_io_warp_ready[1]; // @[pipe.scala 121:59]
  assign ibuffer_io_out_2_ready = ibuffer2issue_io_in_2_ready & warp_sche_io_warp_ready[2]; // @[pipe.scala 121:59]
  assign ibuffer_io_out_3_ready = ibuffer2issue_io_in_3_ready & warp_sche_io_warp_ready[3]; // @[pipe.scala 121:59]
  assign ibuffer2issue_clock = clock;
  assign ibuffer2issue_io_in_0_valid = ibuffer_io_out_0_valid & warp_sche_io_warp_ready[0]; // @[pipe.scala 120:59]
  assign ibuffer2issue_io_in_0_bits_inst = ibuffer_io_out_0_bits_inst; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_wid = ibuffer_io_out_0_bits_wid; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_fp = ibuffer_io_out_0_bits_fp; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_branch = ibuffer_io_out_0_bits_branch; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_simt_stack = ibuffer_io_out_0_bits_simt_stack; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_simt_stack_op = ibuffer_io_out_0_bits_simt_stack_op; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_barrier = ibuffer_io_out_0_bits_barrier; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_csr = ibuffer_io_out_0_bits_csr; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_reverse = ibuffer_io_out_0_bits_reverse; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_sel_alu2 = ibuffer_io_out_0_bits_sel_alu2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_sel_alu1 = ibuffer_io_out_0_bits_sel_alu1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_isvec = ibuffer_io_out_0_bits_isvec; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_sel_alu3 = ibuffer_io_out_0_bits_sel_alu3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_mask = ibuffer_io_out_0_bits_mask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_sel_imm = ibuffer_io_out_0_bits_sel_imm; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_mem_unsigned = ibuffer_io_out_0_bits_mem_unsigned; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_alu_fn = ibuffer_io_out_0_bits_alu_fn; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_mem = ibuffer_io_out_0_bits_mem; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_mem_cmd = ibuffer_io_out_0_bits_mem_cmd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_mop = ibuffer_io_out_0_bits_mop; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_reg_idx1 = ibuffer_io_out_0_bits_reg_idx1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_reg_idx2 = ibuffer_io_out_0_bits_reg_idx2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_reg_idx3 = ibuffer_io_out_0_bits_reg_idx3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_reg_idxw = ibuffer_io_out_0_bits_reg_idxw; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_wfd = ibuffer_io_out_0_bits_wfd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_fence = ibuffer_io_out_0_bits_fence; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_sfu = ibuffer_io_out_0_bits_sfu; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_readmask = ibuffer_io_out_0_bits_readmask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_writemask = ibuffer_io_out_0_bits_writemask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_wxd = ibuffer_io_out_0_bits_wxd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_0_bits_pc = ibuffer_io_out_0_bits_pc; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_valid = ibuffer_io_out_1_valid & warp_sche_io_warp_ready[1]; // @[pipe.scala 120:59]
  assign ibuffer2issue_io_in_1_bits_inst = ibuffer_io_out_1_bits_inst; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_wid = ibuffer_io_out_1_bits_wid; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_fp = ibuffer_io_out_1_bits_fp; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_branch = ibuffer_io_out_1_bits_branch; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_simt_stack = ibuffer_io_out_1_bits_simt_stack; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_simt_stack_op = ibuffer_io_out_1_bits_simt_stack_op; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_barrier = ibuffer_io_out_1_bits_barrier; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_csr = ibuffer_io_out_1_bits_csr; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_reverse = ibuffer_io_out_1_bits_reverse; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_sel_alu2 = ibuffer_io_out_1_bits_sel_alu2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_sel_alu1 = ibuffer_io_out_1_bits_sel_alu1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_isvec = ibuffer_io_out_1_bits_isvec; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_sel_alu3 = ibuffer_io_out_1_bits_sel_alu3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_mask = ibuffer_io_out_1_bits_mask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_sel_imm = ibuffer_io_out_1_bits_sel_imm; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_mem_unsigned = ibuffer_io_out_1_bits_mem_unsigned; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_alu_fn = ibuffer_io_out_1_bits_alu_fn; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_mem = ibuffer_io_out_1_bits_mem; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_mem_cmd = ibuffer_io_out_1_bits_mem_cmd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_mop = ibuffer_io_out_1_bits_mop; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_reg_idx1 = ibuffer_io_out_1_bits_reg_idx1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_reg_idx2 = ibuffer_io_out_1_bits_reg_idx2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_reg_idx3 = ibuffer_io_out_1_bits_reg_idx3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_reg_idxw = ibuffer_io_out_1_bits_reg_idxw; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_wfd = ibuffer_io_out_1_bits_wfd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_fence = ibuffer_io_out_1_bits_fence; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_sfu = ibuffer_io_out_1_bits_sfu; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_readmask = ibuffer_io_out_1_bits_readmask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_writemask = ibuffer_io_out_1_bits_writemask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_wxd = ibuffer_io_out_1_bits_wxd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_1_bits_pc = ibuffer_io_out_1_bits_pc; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_valid = ibuffer_io_out_2_valid & warp_sche_io_warp_ready[2]; // @[pipe.scala 120:59]
  assign ibuffer2issue_io_in_2_bits_inst = ibuffer_io_out_2_bits_inst; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_wid = ibuffer_io_out_2_bits_wid; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_fp = ibuffer_io_out_2_bits_fp; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_branch = ibuffer_io_out_2_bits_branch; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_simt_stack = ibuffer_io_out_2_bits_simt_stack; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_simt_stack_op = ibuffer_io_out_2_bits_simt_stack_op; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_barrier = ibuffer_io_out_2_bits_barrier; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_csr = ibuffer_io_out_2_bits_csr; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_reverse = ibuffer_io_out_2_bits_reverse; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_sel_alu2 = ibuffer_io_out_2_bits_sel_alu2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_sel_alu1 = ibuffer_io_out_2_bits_sel_alu1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_isvec = ibuffer_io_out_2_bits_isvec; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_sel_alu3 = ibuffer_io_out_2_bits_sel_alu3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_mask = ibuffer_io_out_2_bits_mask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_sel_imm = ibuffer_io_out_2_bits_sel_imm; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_mem_unsigned = ibuffer_io_out_2_bits_mem_unsigned; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_alu_fn = ibuffer_io_out_2_bits_alu_fn; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_mem = ibuffer_io_out_2_bits_mem; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_mem_cmd = ibuffer_io_out_2_bits_mem_cmd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_mop = ibuffer_io_out_2_bits_mop; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_reg_idx1 = ibuffer_io_out_2_bits_reg_idx1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_reg_idx2 = ibuffer_io_out_2_bits_reg_idx2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_reg_idx3 = ibuffer_io_out_2_bits_reg_idx3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_reg_idxw = ibuffer_io_out_2_bits_reg_idxw; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_wfd = ibuffer_io_out_2_bits_wfd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_fence = ibuffer_io_out_2_bits_fence; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_sfu = ibuffer_io_out_2_bits_sfu; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_readmask = ibuffer_io_out_2_bits_readmask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_writemask = ibuffer_io_out_2_bits_writemask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_wxd = ibuffer_io_out_2_bits_wxd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_2_bits_pc = ibuffer_io_out_2_bits_pc; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_valid = ibuffer_io_out_3_valid & warp_sche_io_warp_ready[3]; // @[pipe.scala 120:59]
  assign ibuffer2issue_io_in_3_bits_inst = ibuffer_io_out_3_bits_inst; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_wid = ibuffer_io_out_3_bits_wid; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_fp = ibuffer_io_out_3_bits_fp; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_branch = ibuffer_io_out_3_bits_branch; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_simt_stack = ibuffer_io_out_3_bits_simt_stack; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_simt_stack_op = ibuffer_io_out_3_bits_simt_stack_op; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_barrier = ibuffer_io_out_3_bits_barrier; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_csr = ibuffer_io_out_3_bits_csr; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_reverse = ibuffer_io_out_3_bits_reverse; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_sel_alu2 = ibuffer_io_out_3_bits_sel_alu2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_sel_alu1 = ibuffer_io_out_3_bits_sel_alu1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_isvec = ibuffer_io_out_3_bits_isvec; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_sel_alu3 = ibuffer_io_out_3_bits_sel_alu3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_mask = ibuffer_io_out_3_bits_mask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_sel_imm = ibuffer_io_out_3_bits_sel_imm; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_mem_unsigned = ibuffer_io_out_3_bits_mem_unsigned; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_alu_fn = ibuffer_io_out_3_bits_alu_fn; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_mem = ibuffer_io_out_3_bits_mem; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_mem_cmd = ibuffer_io_out_3_bits_mem_cmd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_mop = ibuffer_io_out_3_bits_mop; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_reg_idx1 = ibuffer_io_out_3_bits_reg_idx1; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_reg_idx2 = ibuffer_io_out_3_bits_reg_idx2; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_reg_idx3 = ibuffer_io_out_3_bits_reg_idx3; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_reg_idxw = ibuffer_io_out_3_bits_reg_idxw; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_wfd = ibuffer_io_out_3_bits_wfd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_fence = ibuffer_io_out_3_bits_fence; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_sfu = ibuffer_io_out_3_bits_sfu; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_readmask = ibuffer_io_out_3_bits_readmask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_writemask = ibuffer_io_out_3_bits_writemask; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_wxd = ibuffer_io_out_3_bits_wxd; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_in_3_bits_pc = ibuffer_io_out_3_bits_pc; // @[pipe.scala 119:32]
  assign ibuffer2issue_io_out_ready = exe_data_io_enq_ready; // @[pipe.scala 213:29]
  assign exe_data_clock = clock;
  assign exe_data_reset = reset;
  assign exe_data_io_enq_valid = ibuffer2issue_io_out_valid; // @[pipe.scala 211:26]
  assign exe_data_io_enq_bits_in1_0 = operand_collector_io_alu_src1_0; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_1 = operand_collector_io_alu_src1_1; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_2 = operand_collector_io_alu_src1_2; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_3 = operand_collector_io_alu_src1_3; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_4 = operand_collector_io_alu_src1_4; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_5 = operand_collector_io_alu_src1_5; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_6 = operand_collector_io_alu_src1_6; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in1_7 = operand_collector_io_alu_src1_7; // @[pipe.scala 207:30]
  assign exe_data_io_enq_bits_in2_0 = operand_collector_io_alu_src2_0; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_1 = operand_collector_io_alu_src2_1; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_2 = operand_collector_io_alu_src2_2; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_3 = operand_collector_io_alu_src2_3; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_4 = operand_collector_io_alu_src2_4; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_5 = operand_collector_io_alu_src2_5; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_6 = operand_collector_io_alu_src2_6; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in2_7 = operand_collector_io_alu_src2_7; // @[pipe.scala 208:30]
  assign exe_data_io_enq_bits_in3_0 = operand_collector_io_alu_src3_0; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_1 = operand_collector_io_alu_src3_1; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_2 = operand_collector_io_alu_src3_2; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_3 = operand_collector_io_alu_src3_3; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_4 = operand_collector_io_alu_src3_4; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_5 = operand_collector_io_alu_src3_5; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_6 = operand_collector_io_alu_src3_6; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_in3_7 = operand_collector_io_alu_src3_7; // @[pipe.scala 209:30]
  assign exe_data_io_enq_bits_mask_0 = operand_collector_io_mask_0 & simt_stack_io_out_mask[0]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_1 = operand_collector_io_mask_1 & simt_stack_io_out_mask[1]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_2 = operand_collector_io_mask_2 & simt_stack_io_out_mask[2]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_3 = operand_collector_io_mask_3 & simt_stack_io_out_mask[3]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_4 = operand_collector_io_mask_4 & simt_stack_io_out_mask[4]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_5 = operand_collector_io_mask_5 & simt_stack_io_out_mask[5]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_6 = operand_collector_io_mask_6 & simt_stack_io_out_mask[6]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_mask_7 = operand_collector_io_mask_7 & simt_stack_io_out_mask[7]; // @[pipe.scala 210:90]
  assign exe_data_io_enq_bits_ctrl_inst = ibuffer2issue_io_out_bits_inst; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_wid = ibuffer2issue_io_out_bits_wid; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_fp = ibuffer2issue_io_out_bits_fp; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_branch = ibuffer2issue_io_out_bits_branch; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_simt_stack = ibuffer2issue_io_out_bits_simt_stack; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_simt_stack_op = ibuffer2issue_io_out_bits_simt_stack_op; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_barrier = ibuffer2issue_io_out_bits_barrier; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_csr = ibuffer2issue_io_out_bits_csr; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_reverse = ibuffer2issue_io_out_bits_reverse; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_isvec = ibuffer2issue_io_out_bits_isvec; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_mem_unsigned = ibuffer2issue_io_out_bits_mem_unsigned; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_alu_fn = ibuffer2issue_io_out_bits_alu_fn; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_mem = ibuffer2issue_io_out_bits_mem; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_mem_cmd = ibuffer2issue_io_out_bits_mem_cmd; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_mop = ibuffer2issue_io_out_bits_mop; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_reg_idxw = ibuffer2issue_io_out_bits_reg_idxw; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_wfd = ibuffer2issue_io_out_bits_wfd; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_fence = ibuffer2issue_io_out_bits_fence; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_sfu = ibuffer2issue_io_out_bits_sfu; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_readmask = ibuffer2issue_io_out_bits_readmask; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_writemask = ibuffer2issue_io_out_bits_writemask; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_wxd = ibuffer2issue_io_out_bits_wxd; // @[pipe.scala 206:31]
  assign exe_data_io_enq_bits_ctrl_pc = ibuffer2issue_io_out_bits_pc; // @[pipe.scala 206:31]
  assign exe_data_io_deq_ready = issue_io_in_ready; // @[pipe.scala 214:14]
  assign simt_stack_clock = clock;
  assign simt_stack_reset = reset;
  assign simt_stack_io_branch_ctl_valid = issue_io_out_SIMT_valid; // @[pipe.scala 220:20]
  assign simt_stack_io_branch_ctl_bits_opcode = issue_io_out_SIMT_bits_opcode; // @[pipe.scala 220:20]
  assign simt_stack_io_branch_ctl_bits_wid = issue_io_out_SIMT_bits_wid; // @[pipe.scala 220:20]
  assign simt_stack_io_branch_ctl_bits_PC_branch = issue_io_out_SIMT_bits_PC_branch; // @[pipe.scala 220:20]
  assign simt_stack_io_branch_ctl_bits_mask_init = issue_io_out_SIMT_bits_mask_init; // @[pipe.scala 220:20]
  assign simt_stack_io_if_mask_valid = valu_io_out2simt_stack_valid; // @[pipe.scala 223:24]
  assign simt_stack_io_if_mask_bits_if_mask = valu_io_out2simt_stack_bits_if_mask; // @[pipe.scala 223:24]
  assign simt_stack_io_if_mask_bits_wid = valu_io_out2simt_stack_bits_wid; // @[pipe.scala 223:24]
  assign simt_stack_io_input_wid = ibuffer2issue_io_out_bits_wid; // @[pipe.scala 155:26]
  assign simt_stack_io_fetch_ctl_ready = branch_back_io_in1_ready; // @[pipe.scala 224:26]
  assign branch_back_io_out_ready = warp_sche_io_branch_ready; // @[pipe.scala 64:22]
  assign branch_back_io_in0_valid = alu_io_out2br_valid; // @[pipe.scala 226:16]
  assign branch_back_io_in0_bits_wid = alu_io_out2br_bits_wid; // @[pipe.scala 226:16]
  assign branch_back_io_in0_bits_jump = alu_io_out2br_bits_jump; // @[pipe.scala 226:16]
  assign branch_back_io_in0_bits_new_pc = alu_io_out2br_bits_new_pc; // @[pipe.scala 226:16]
  assign branch_back_io_in1_valid = simt_stack_io_fetch_ctl_valid; // @[pipe.scala 224:26]
  assign branch_back_io_in1_bits_wid = simt_stack_io_fetch_ctl_bits_wid; // @[pipe.scala 224:26]
  assign branch_back_io_in1_bits_jump = simt_stack_io_fetch_ctl_bits_jump; // @[pipe.scala 224:26]
  assign branch_back_io_in1_bits_new_pc = simt_stack_io_fetch_ctl_bits_new_pc; // @[pipe.scala 224:26]
  assign csrfile_clock = clock;
  assign csrfile_reset = reset;
  assign csrfile_io_in_valid = issue_io_out_CSR_valid; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_ctrl_inst = issue_io_out_CSR_bits_ctrl_inst; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_ctrl_wid = issue_io_out_CSR_bits_ctrl_wid; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_ctrl_csr = issue_io_out_CSR_bits_ctrl_csr; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_ctrl_isvec = issue_io_out_CSR_bits_ctrl_isvec; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_ctrl_reg_idxw = issue_io_out_CSR_bits_ctrl_reg_idxw; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_ctrl_wxd = issue_io_out_CSR_bits_ctrl_wxd; // @[pipe.scala 219:19]
  assign csrfile_io_in_bits_in1 = issue_io_out_CSR_bits_in1; // @[pipe.scala 219:19]
  assign csrfile_io_out_ready = wb_io_in_x_3_ready; // @[pipe.scala 242:16]
  assign csrfile_io_frm_wid = fpu_io_in_bits_ctrl_wid; // @[pipe.scala 231:21]
  assign csrfile_io_CTA2csr_valid = warp_sche_io_CTA2csr_valid; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count =
    warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wg_wf_count; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    warp_sche_io_CTA2csr_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[pipe.scala 79:21]
  assign csrfile_io_CTA2csr_bits_wid = warp_sche_io_CTA2csr_bits_wid; // @[pipe.scala 79:21]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset) begin
          $fwrite(32'h80000002,"undefined instructions at 0x%x with 0x%x\n",control_io_pc,control_io_inst); // @[pipe.scala 102:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"0x%x,writedata=",exe_data_io_deq_bits_ctrl_pc); // @[pipe.scala 187:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_0); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_1); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_2); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_3); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_4); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_5); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_6); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in2_7); // @[pipe.scala 188:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_0); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_1); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_2); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_3); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_4); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_5); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_6); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in1_7); // @[pipe.scala 189:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_0); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_1); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_2); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_3); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_4); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_5); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_6); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_in3_7); // @[pipe.scala 190:48]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_0); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_1); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_2); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_3); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_4); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_5); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_6); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"%x ",exe_data_io_deq_bits_mask_7); // @[pipe.scala 191:49]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_3) begin
          $fwrite(32'h80000002,"\n"); // @[pipe.scala 192:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter_14(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_a_addr,
  input  [2:0]  io_in_0_bits_a_source,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [2:0]  io_in_1_bits_a_opcode,
  input  [31:0] io_in_1_bits_a_addr,
  input  [31:0] io_in_1_bits_a_data_0,
  input  [31:0] io_in_1_bits_a_data_1,
  input  [31:0] io_in_1_bits_a_data_2,
  input  [31:0] io_in_1_bits_a_data_3,
  input  [31:0] io_in_1_bits_a_data_4,
  input  [31:0] io_in_1_bits_a_data_5,
  input  [31:0] io_in_1_bits_a_data_6,
  input  [31:0] io_in_1_bits_a_data_7,
  input         io_in_1_bits_a_mask_0,
  input         io_in_1_bits_a_mask_1,
  input         io_in_1_bits_a_mask_2,
  input         io_in_1_bits_a_mask_3,
  input         io_in_1_bits_a_mask_4,
  input         io_in_1_bits_a_mask_5,
  input         io_in_1_bits_a_mask_6,
  input         io_in_1_bits_a_mask_7,
  input  [2:0]  io_in_1_bits_a_source,
  input         io_out_ready,
  output        io_out_valid,
  output [2:0]  io_out_bits_a_opcode,
  output [31:0] io_out_bits_a_addr,
  output [31:0] io_out_bits_a_data_0,
  output [31:0] io_out_bits_a_data_1,
  output [31:0] io_out_bits_a_data_2,
  output [31:0] io_out_bits_a_data_3,
  output [31:0] io_out_bits_a_data_4,
  output [31:0] io_out_bits_a_data_5,
  output [31:0] io_out_bits_a_data_6,
  output [31:0] io_out_bits_a_data_7,
  output        io_out_bits_a_mask_0,
  output        io_out_bits_a_mask_1,
  output        io_out_bits_a_mask_2,
  output        io_out_bits_a_mask_3,
  output        io_out_bits_a_mask_4,
  output        io_out_bits_a_mask_5,
  output        io_out_bits_a_mask_6,
  output        io_out_bits_a_mask_7,
  output [2:0]  io_out_bits_a_source
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_a_opcode = io_in_0_valid ? 3'h4 : io_in_1_bits_a_opcode; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_addr = io_in_0_valid ? io_in_0_bits_a_addr : io_in_1_bits_a_addr; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_0 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_0; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_1 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_1; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_2 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_2; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_3 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_3; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_4 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_4; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_5 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_5; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_6 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_6; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_7 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_7; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_0 = io_in_0_valid | io_in_1_bits_a_mask_0; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_1 = io_in_0_valid | io_in_1_bits_a_mask_1; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_2 = io_in_0_valid | io_in_1_bits_a_mask_2; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_3 = io_in_0_valid | io_in_1_bits_a_mask_3; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_4 = io_in_0_valid | io_in_1_bits_a_mask_4; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_5 = io_in_0_valid | io_in_1_bits_a_mask_5; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_6 = io_in_0_valid | io_in_1_bits_a_mask_6; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_7 = io_in_0_valid | io_in_1_bits_a_mask_7; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_source = io_in_0_valid ? io_in_0_bits_a_source : io_in_1_bits_a_source; // @[Arbiter.scala 139:15 141:26 143:19]
endmodule
module L1Cache2L2Arbiter(
  output        io_memReqVecIn_0_ready,
  input         io_memReqVecIn_0_valid,
  input  [1:0]  io_memReqVecIn_0_bits_a_source,
  input  [31:0] io_memReqVecIn_0_bits_a_addr,
  output        io_memReqVecIn_1_ready,
  input         io_memReqVecIn_1_valid,
  input  [2:0]  io_memReqVecIn_1_bits_a_opcode,
  input  [1:0]  io_memReqVecIn_1_bits_a_source,
  input  [31:0] io_memReqVecIn_1_bits_a_addr,
  input  [31:0] io_memReqVecIn_1_bits_a_data_0,
  input  [31:0] io_memReqVecIn_1_bits_a_data_1,
  input  [31:0] io_memReqVecIn_1_bits_a_data_2,
  input  [31:0] io_memReqVecIn_1_bits_a_data_3,
  input  [31:0] io_memReqVecIn_1_bits_a_data_4,
  input  [31:0] io_memReqVecIn_1_bits_a_data_5,
  input  [31:0] io_memReqVecIn_1_bits_a_data_6,
  input  [31:0] io_memReqVecIn_1_bits_a_data_7,
  input         io_memReqVecIn_1_bits_a_mask_0,
  input         io_memReqVecIn_1_bits_a_mask_1,
  input         io_memReqVecIn_1_bits_a_mask_2,
  input         io_memReqVecIn_1_bits_a_mask_3,
  input         io_memReqVecIn_1_bits_a_mask_4,
  input         io_memReqVecIn_1_bits_a_mask_5,
  input         io_memReqVecIn_1_bits_a_mask_6,
  input         io_memReqVecIn_1_bits_a_mask_7,
  input         io_memReqOut_ready,
  output        io_memReqOut_valid,
  output [2:0]  io_memReqOut_bits_a_opcode,
  output [31:0] io_memReqOut_bits_a_addr,
  output [31:0] io_memReqOut_bits_a_data_0,
  output [31:0] io_memReqOut_bits_a_data_1,
  output [31:0] io_memReqOut_bits_a_data_2,
  output [31:0] io_memReqOut_bits_a_data_3,
  output [31:0] io_memReqOut_bits_a_data_4,
  output [31:0] io_memReqOut_bits_a_data_5,
  output [31:0] io_memReqOut_bits_a_data_6,
  output [31:0] io_memReqOut_bits_a_data_7,
  output        io_memReqOut_bits_a_mask_0,
  output        io_memReqOut_bits_a_mask_1,
  output        io_memReqOut_bits_a_mask_2,
  output        io_memReqOut_bits_a_mask_3,
  output        io_memReqOut_bits_a_mask_4,
  output        io_memReqOut_bits_a_mask_5,
  output        io_memReqOut_bits_a_mask_6,
  output        io_memReqOut_bits_a_mask_7,
  output [2:0]  io_memReqOut_bits_a_source,
  output        io_memRspIn_ready,
  input         io_memRspIn_valid,
  input  [31:0] io_memRspIn_bits_d_addr,
  input  [31:0] io_memRspIn_bits_d_data_0,
  input  [31:0] io_memRspIn_bits_d_data_1,
  input  [31:0] io_memRspIn_bits_d_data_2,
  input  [31:0] io_memRspIn_bits_d_data_3,
  input  [31:0] io_memRspIn_bits_d_data_4,
  input  [31:0] io_memRspIn_bits_d_data_5,
  input  [31:0] io_memRspIn_bits_d_data_6,
  input  [31:0] io_memRspIn_bits_d_data_7,
  input  [2:0]  io_memRspIn_bits_d_source,
  input         io_memRspVecOut_0_ready,
  output        io_memRspVecOut_0_valid,
  output [31:0] io_memRspVecOut_0_bits_d_addr,
  output [31:0] io_memRspVecOut_0_bits_d_data_0,
  output [31:0] io_memRspVecOut_0_bits_d_data_1,
  output [31:0] io_memRspVecOut_0_bits_d_data_2,
  output [31:0] io_memRspVecOut_0_bits_d_data_3,
  output [31:0] io_memRspVecOut_0_bits_d_data_4,
  output [31:0] io_memRspVecOut_0_bits_d_data_5,
  output [31:0] io_memRspVecOut_0_bits_d_data_6,
  output [31:0] io_memRspVecOut_0_bits_d_data_7,
  input         io_memRspVecOut_1_ready,
  output        io_memRspVecOut_1_valid,
  output [31:0] io_memRspVecOut_1_bits_d_addr,
  output [31:0] io_memRspVecOut_1_bits_d_data_0,
  output [31:0] io_memRspVecOut_1_bits_d_data_1,
  output [31:0] io_memRspVecOut_1_bits_d_data_2,
  output [31:0] io_memRspVecOut_1_bits_d_data_3,
  output [31:0] io_memRspVecOut_1_bits_d_data_4,
  output [31:0] io_memRspVecOut_1_bits_d_data_5,
  output [31:0] io_memRspVecOut_1_bits_d_data_6,
  output [31:0] io_memRspVecOut_1_bits_d_data_7
);
  wire  memReqArb_io_in_0_ready; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_0_valid; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_0_bits_a_addr; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [2:0] memReqArb_io_in_0_bits_a_source; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_ready; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_valid; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [2:0] memReqArb_io_in_1_bits_a_opcode; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_addr; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_0; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_1; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_2; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_3; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_4; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_5; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_6; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_in_1_bits_a_data_7; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_0; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_1; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_2; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_3; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_4; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_5; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_6; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_in_1_bits_a_mask_7; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [2:0] memReqArb_io_in_1_bits_a_source; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_ready; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_valid; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [2:0] memReqArb_io_out_bits_a_opcode; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_addr; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_0; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_1; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_2; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_3; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_4; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_5; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_6; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [31:0] memReqArb_io_out_bits_a_data_7; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_0; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_1; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_2; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_3; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_4; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_5; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_6; // @[L1Cache2L2Arbiter.scala 27:25]
  wire  memReqArb_io_out_bits_a_mask_7; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [2:0] memReqArb_io_out_bits_a_source; // @[L1Cache2L2Arbiter.scala 27:25]
  wire [1:0] _io_memRspIn_ready_T_1 = 2'h1 << io_memRspIn_bits_d_source[2]; // @[OneHot.scala 57:35]
  wire [1:0] _io_memRspIn_ready_T_2 = {io_memRspVecOut_0_ready,io_memRspVecOut_1_ready}; // @[Cat.scala 31:58]
  wire [1:0] _io_memRspIn_ready_T_5 = {_io_memRspIn_ready_T_2[0],_io_memRspIn_ready_T_2[1]}; // @[Cat.scala 31:58]
  wire [1:0] _io_memRspIn_ready_T_6 = _io_memRspIn_ready_T_1 & _io_memRspIn_ready_T_5; // @[Mux.scala 30:47]
  Arbiter_14 memReqArb ( // @[L1Cache2L2Arbiter.scala 27:25]
    .io_in_0_ready(memReqArb_io_in_0_ready),
    .io_in_0_valid(memReqArb_io_in_0_valid),
    .io_in_0_bits_a_addr(memReqArb_io_in_0_bits_a_addr),
    .io_in_0_bits_a_source(memReqArb_io_in_0_bits_a_source),
    .io_in_1_ready(memReqArb_io_in_1_ready),
    .io_in_1_valid(memReqArb_io_in_1_valid),
    .io_in_1_bits_a_opcode(memReqArb_io_in_1_bits_a_opcode),
    .io_in_1_bits_a_addr(memReqArb_io_in_1_bits_a_addr),
    .io_in_1_bits_a_data_0(memReqArb_io_in_1_bits_a_data_0),
    .io_in_1_bits_a_data_1(memReqArb_io_in_1_bits_a_data_1),
    .io_in_1_bits_a_data_2(memReqArb_io_in_1_bits_a_data_2),
    .io_in_1_bits_a_data_3(memReqArb_io_in_1_bits_a_data_3),
    .io_in_1_bits_a_data_4(memReqArb_io_in_1_bits_a_data_4),
    .io_in_1_bits_a_data_5(memReqArb_io_in_1_bits_a_data_5),
    .io_in_1_bits_a_data_6(memReqArb_io_in_1_bits_a_data_6),
    .io_in_1_bits_a_data_7(memReqArb_io_in_1_bits_a_data_7),
    .io_in_1_bits_a_mask_0(memReqArb_io_in_1_bits_a_mask_0),
    .io_in_1_bits_a_mask_1(memReqArb_io_in_1_bits_a_mask_1),
    .io_in_1_bits_a_mask_2(memReqArb_io_in_1_bits_a_mask_2),
    .io_in_1_bits_a_mask_3(memReqArb_io_in_1_bits_a_mask_3),
    .io_in_1_bits_a_mask_4(memReqArb_io_in_1_bits_a_mask_4),
    .io_in_1_bits_a_mask_5(memReqArb_io_in_1_bits_a_mask_5),
    .io_in_1_bits_a_mask_6(memReqArb_io_in_1_bits_a_mask_6),
    .io_in_1_bits_a_mask_7(memReqArb_io_in_1_bits_a_mask_7),
    .io_in_1_bits_a_source(memReqArb_io_in_1_bits_a_source),
    .io_out_ready(memReqArb_io_out_ready),
    .io_out_valid(memReqArb_io_out_valid),
    .io_out_bits_a_opcode(memReqArb_io_out_bits_a_opcode),
    .io_out_bits_a_addr(memReqArb_io_out_bits_a_addr),
    .io_out_bits_a_data_0(memReqArb_io_out_bits_a_data_0),
    .io_out_bits_a_data_1(memReqArb_io_out_bits_a_data_1),
    .io_out_bits_a_data_2(memReqArb_io_out_bits_a_data_2),
    .io_out_bits_a_data_3(memReqArb_io_out_bits_a_data_3),
    .io_out_bits_a_data_4(memReqArb_io_out_bits_a_data_4),
    .io_out_bits_a_data_5(memReqArb_io_out_bits_a_data_5),
    .io_out_bits_a_data_6(memReqArb_io_out_bits_a_data_6),
    .io_out_bits_a_data_7(memReqArb_io_out_bits_a_data_7),
    .io_out_bits_a_mask_0(memReqArb_io_out_bits_a_mask_0),
    .io_out_bits_a_mask_1(memReqArb_io_out_bits_a_mask_1),
    .io_out_bits_a_mask_2(memReqArb_io_out_bits_a_mask_2),
    .io_out_bits_a_mask_3(memReqArb_io_out_bits_a_mask_3),
    .io_out_bits_a_mask_4(memReqArb_io_out_bits_a_mask_4),
    .io_out_bits_a_mask_5(memReqArb_io_out_bits_a_mask_5),
    .io_out_bits_a_mask_6(memReqArb_io_out_bits_a_mask_6),
    .io_out_bits_a_mask_7(memReqArb_io_out_bits_a_mask_7),
    .io_out_bits_a_source(memReqArb_io_out_bits_a_source)
  );
  assign io_memReqVecIn_0_ready = memReqArb_io_in_0_ready; // @[L1Cache2L2Arbiter.scala 28:19]
  assign io_memReqVecIn_1_ready = memReqArb_io_in_1_ready; // @[L1Cache2L2Arbiter.scala 28:19]
  assign io_memReqOut_valid = memReqArb_io_out_valid; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_opcode = memReqArb_io_out_bits_a_opcode; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_addr = memReqArb_io_out_bits_a_addr; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_0 = memReqArb_io_out_bits_a_data_0; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_1 = memReqArb_io_out_bits_a_data_1; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_2 = memReqArb_io_out_bits_a_data_2; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_3 = memReqArb_io_out_bits_a_data_3; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_4 = memReqArb_io_out_bits_a_data_4; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_5 = memReqArb_io_out_bits_a_data_5; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_6 = memReqArb_io_out_bits_a_data_6; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_data_7 = memReqArb_io_out_bits_a_data_7; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_0 = memReqArb_io_out_bits_a_mask_0; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_1 = memReqArb_io_out_bits_a_mask_1; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_2 = memReqArb_io_out_bits_a_mask_2; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_3 = memReqArb_io_out_bits_a_mask_3; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_4 = memReqArb_io_out_bits_a_mask_4; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_5 = memReqArb_io_out_bits_a_mask_5; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_6 = memReqArb_io_out_bits_a_mask_6; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_mask_7 = memReqArb_io_out_bits_a_mask_7; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memReqOut_bits_a_source = memReqArb_io_out_bits_a_source; // @[L1Cache2L2Arbiter.scala 32:16]
  assign io_memRspIn_ready = |_io_memRspIn_ready_T_6; // @[Mux.scala 30:53]
  assign io_memRspVecOut_0_valid = ~io_memRspIn_bits_d_source[2] & io_memRspIn_valid; // @[L1Cache2L2Arbiter.scala 39:82]
  assign io_memRspVecOut_0_bits_d_addr = io_memRspIn_bits_d_addr; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_0 = io_memRspIn_bits_d_data_0; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_1 = io_memRspIn_bits_d_data_1; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_2 = io_memRspIn_bits_d_data_2; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_3 = io_memRspIn_bits_d_data_3; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_4 = io_memRspIn_bits_d_data_4; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_5 = io_memRspIn_bits_d_data_5; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_6 = io_memRspIn_bits_d_data_6; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_0_bits_d_data_7 = io_memRspIn_bits_d_data_7; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_valid = io_memRspIn_bits_d_source[2] & io_memRspIn_valid; // @[L1Cache2L2Arbiter.scala 39:82]
  assign io_memRspVecOut_1_bits_d_addr = io_memRspIn_bits_d_addr; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_0 = io_memRspIn_bits_d_data_0; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_1 = io_memRspIn_bits_d_data_1; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_2 = io_memRspIn_bits_d_data_2; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_3 = io_memRspIn_bits_d_data_3; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_4 = io_memRspIn_bits_d_data_4; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_5 = io_memRspIn_bits_d_data_5; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_6 = io_memRspIn_bits_d_data_6; // @[L1Cache2L2Arbiter.scala 37:29]
  assign io_memRspVecOut_1_bits_d_data_7 = io_memRspIn_bits_d_data_7; // @[L1Cache2L2Arbiter.scala 37:29]
  assign memReqArb_io_in_0_valid = io_memReqVecIn_0_valid; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_0_bits_a_addr = io_memReqVecIn_0_bits_a_addr; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_0_bits_a_source = {1'h0,io_memReqVecIn_0_bits_a_source}; // @[Cat.scala 31:58]
  assign memReqArb_io_in_1_valid = io_memReqVecIn_1_valid; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_opcode = io_memReqVecIn_1_bits_a_opcode; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_addr = io_memReqVecIn_1_bits_a_addr; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_0 = io_memReqVecIn_1_bits_a_data_0; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_1 = io_memReqVecIn_1_bits_a_data_1; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_2 = io_memReqVecIn_1_bits_a_data_2; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_3 = io_memReqVecIn_1_bits_a_data_3; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_4 = io_memReqVecIn_1_bits_a_data_4; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_5 = io_memReqVecIn_1_bits_a_data_5; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_6 = io_memReqVecIn_1_bits_a_data_6; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_data_7 = io_memReqVecIn_1_bits_a_data_7; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_0 = io_memReqVecIn_1_bits_a_mask_0; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_1 = io_memReqVecIn_1_bits_a_mask_1; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_2 = io_memReqVecIn_1_bits_a_mask_2; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_3 = io_memReqVecIn_1_bits_a_mask_3; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_4 = io_memReqVecIn_1_bits_a_mask_4; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_5 = io_memReqVecIn_1_bits_a_mask_5; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_6 = io_memReqVecIn_1_bits_a_mask_6; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_mask_7 = io_memReqVecIn_1_bits_a_mask_7; // @[L1Cache2L2Arbiter.scala 28:19]
  assign memReqArb_io_in_1_bits_a_source = {1'h1,io_memReqVecIn_1_bits_a_source}; // @[Cat.scala 31:58]
  assign memReqArb_io_out_ready = io_memReqOut_ready; // @[L1Cache2L2Arbiter.scala 32:16]
endmodule
module SRAMTemplate(
  input         clock,
  input         reset,
  input         io_r_req_valid,
  input  [4:0]  io_r_req_bits_setIdx,
  output [21:0] io_r_resp_data_0,
  output [21:0] io_r_resp_data_1,
  input         io_w_req_valid,
  input  [4:0]  io_w_req_bits_setIdx,
  input  [21:0] io_w_req_bits_data_0,
  input  [21:0] io_w_req_bits_data_1,
  input  [1:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] array_0 [0:31]; // @[SRAMTemplate.scala 101:26]
  wire  array_0_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_0_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [21:0] array_0_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [21:0] array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_0_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_0_raw_rdata_en_pipe_0;
  reg [4:0] array_0_raw_rdata_addr_pipe_0;
  reg [21:0] array_1 [0:31]; // @[SRAMTemplate.scala 101:26]
  wire  array_1_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_1_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [21:0] array_1_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [21:0] array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_1_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_1_raw_rdata_en_pipe_0;
  reg [4:0] array_1_raw_rdata_addr_pipe_0;
  reg [63:0] bypass_wdata_lfsr; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor = bypass_wdata_lfsr[0] ^ bypass_wdata_lfsr[1] ^ bypass_wdata_lfsr[3] ^ bypass_wdata_lfsr[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_2 = {bypass_wdata_xor,bypass_wdata_lfsr[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_1; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_1 = bypass_wdata_lfsr_1[0] ^ bypass_wdata_lfsr_1[1] ^ bypass_wdata_lfsr_1[3] ^
    bypass_wdata_lfsr_1[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_6 = {bypass_wdata_xor_1,bypass_wdata_lfsr_1[63:1]}; // @[Cat.scala 31:58]
  reg  bypass_mask_need_check; // @[SRAMTemplate.scala 126:29]
  reg [4:0] bypass_mask_waddr_reg; // @[SRAMTemplate.scala 127:28]
  reg [4:0] bypass_mask_raddr_reg; // @[SRAMTemplate.scala 128:28]
  wire  _bypass_mask_bypass_T_1 = bypass_mask_need_check & bypass_mask_waddr_reg == bypass_mask_raddr_reg; // @[SRAMTemplate.scala 130:39]
  wire [1:0] _bypass_mask_bypass_T_3 = _bypass_mask_bypass_T_1 ? 2'h3 : 2'h0; // @[Bitwise.scala 74:12]
  reg [1:0] bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:76]
  wire [1:0] bypass_mask_bypass = _bypass_mask_bypass_T_3 & bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:67]
  wire [21:0] bypass_wdata_0 = bypass_wdata_lfsr[21:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [21:0] mem_rdata_0 = bypass_mask_bypass[0] ? bypass_wdata_0 : array_0_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  wire [21:0] bypass_wdata_1 = bypass_wdata_lfsr_1[21:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [21:0] mem_rdata_1 = bypass_mask_bypass[1] ? bypass_wdata_1 : array_1_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  reg  rdata_REG; // @[SRAMTemplate.scala 144:59]
  reg [21:0] rdata_r_0; // @[Reg.scala 28:20]
  reg [21:0] rdata_r_1; // @[Reg.scala 28:20]
  assign array_0_raw_rdata_en = array_0_raw_rdata_en_pipe_0;
  assign array_0_raw_rdata_addr = array_0_raw_rdata_addr_pipe_0;
  assign array_0_raw_rdata_data = array_0[array_0_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_0_MPORT_data = io_w_req_bits_data_0;
  assign array_0_MPORT_addr = io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = io_w_req_bits_waymask[0];
  assign array_0_MPORT_en = io_w_req_valid;
  assign array_1_raw_rdata_en = array_1_raw_rdata_en_pipe_0;
  assign array_1_raw_rdata_addr = array_1_raw_rdata_addr_pipe_0;
  assign array_1_raw_rdata_data = array_1[array_1_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_1_MPORT_data = io_w_req_bits_data_1;
  assign array_1_MPORT_addr = io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = io_w_req_bits_waymask[1];
  assign array_1_MPORT_en = io_w_req_valid;
  assign io_r_resp_data_0 = rdata_REG ? mem_rdata_0 : rdata_r_0; // @[Hold.scala 23:48]
  assign io_r_resp_data_1 = rdata_REG ? mem_rdata_1 : rdata_r_1; // @[Hold.scala 23:48]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_0_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_0_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_1_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_1_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr <= 64'h1;
    end else begin
      bypass_wdata_lfsr <= _bypass_wdata_lfsr_T_2;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_1 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_1 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_1 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_1 <= _bypass_wdata_lfsr_T_6;
    end
    bypass_mask_need_check <= io_r_req_valid & io_w_req_valid; // @[SRAMTemplate.scala 126:34]
    bypass_mask_waddr_reg <= io_w_req_bits_setIdx; // @[SRAMTemplate.scala 127:28]
    bypass_mask_raddr_reg <= io_r_req_bits_setIdx; // @[SRAMTemplate.scala 128:28]
    bypass_mask_bypass_REG <= io_w_req_bits_waymask; // @[SRAMTemplate.scala 130:76]
    rdata_REG <= io_r_req_valid; // @[SRAMTemplate.scala 144:59]
    if (reset) begin // @[Reg.scala 28:20]
      rdata_r_0 <= 22'h0; // @[Reg.scala 28:20]
    end else if (rdata_REG) begin // @[Reg.scala 29:18]
      if (bypass_mask_bypass[0]) begin // @[SRAMTemplate.scala 139:30]
        rdata_r_0 <= bypass_wdata_0;
      end else begin
        rdata_r_0 <= array_0_raw_rdata_data;
      end
    end
    if (reset) begin // @[Reg.scala 28:20]
      rdata_r_1 <= 22'h0; // @[Reg.scala 28:20]
    end else if (rdata_REG) begin // @[Reg.scala 29:18]
      if (bypass_mask_bypass[1]) begin // @[SRAMTemplate.scala 139:30]
        rdata_r_1 <= bypass_wdata_1;
      end else begin
        rdata_r_1 <= array_1_raw_rdata_data;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    array_0[initvar] = _RAND_0[21:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    array_1[initvar] = _RAND_3[21:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_raw_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_raw_rdata_addr_pipe_0 = _RAND_2[4:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_raw_rdata_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_raw_rdata_addr_pipe_0 = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  bypass_wdata_lfsr = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  bypass_wdata_lfsr_1 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  bypass_mask_need_check = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  bypass_mask_waddr_reg = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  bypass_mask_raddr_reg = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  bypass_mask_bypass_REG = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  rdata_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rdata_r_0 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  rdata_r_1 = _RAND_14[21:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module tagChecker(
  input         clock,
  input         reset,
  input  [21:0] io_tag_of_set_0,
  input  [21:0] io_tag_of_set_1,
  input  [21:0] io_tag_from_pipe,
  input         io_way_valid_0,
  input         io_way_valid_1,
  output [1:0]  io_waymask,
  output        io_cache_hit
);
  wire  _io_waymask_T_1 = io_tag_of_set_0 == io_tag_from_pipe & io_way_valid_0; // @[L1CacheSubModules.scala 98:112]
  wire  _io_waymask_T_3 = io_tag_of_set_1 == io_tag_from_pipe & io_way_valid_1; // @[L1CacheSubModules.scala 98:112]
  wire [1:0] _io_waymask_T_4 = {_io_waymask_T_1,_io_waymask_T_3}; // @[Cat.scala 31:58]
  wire [1:0] _T_2 = io_waymask[0] + io_waymask[1]; // @[Bitwise.scala 48:55]
  assign io_waymask = {_io_waymask_T_4[0],_io_waymask_T_4[1]}; // @[Cat.scala 31:58]
  assign io_cache_hit = |io_waymask; // @[L1CacheSubModules.scala 101:30]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(_T_2 <= 2'h1)) begin
          $fatal; // @[L1CacheSubModules.scala 100:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_2 <= 2'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at L1CacheSubModules.scala:100 assert(PopCount(io.waymask) <= 1.U)//if waymask not one-hot, duplicate tags in one set, error\n"
            ); // @[L1CacheSubModules.scala 100:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ReplacementUnit(
  input        clock,
  input        reset,
  input  [1:0] io_validbits_of_set,
  output [1:0] io_waymask,
  output       io_Set_is_full
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] victim_1Hidx; // @[L1CacheSubModules.scala 79:40]
  wire  _io_waymask_T_4 = ~io_validbits_of_set[0] ? 1'h0 : 1'h1; // @[L1CacheSubModules.scala 81:107]
  wire [1:0] _io_waymask_T_5 = 2'h1 << _io_waymask_T_4; // @[OneHot.scala 57:35]
  wire [1:0] _victim_1Hidx_T_2 = {victim_1Hidx[0],victim_1Hidx[1]}; // @[Cat.scala 31:58]
  reg [1:0] victim_1Hidx_r; // @[Reg.scala 16:16]
  assign io_waymask = io_Set_is_full ? victim_1Hidx : _io_waymask_T_5; // @[L1CacheSubModules.scala 81:20]
  assign io_Set_is_full = io_validbits_of_set == 2'h3; // @[L1CacheSubModules.scala 80:41]
  always @(posedge clock) begin
    if (reset) begin // @[L1CacheSubModules.scala 79:40]
      victim_1Hidx <= 2'h1; // @[L1CacheSubModules.scala 79:40]
    end else begin
      victim_1Hidx <= victim_1Hidx_r; // @[L1CacheSubModules.scala 84:27]
    end
    if (io_Set_is_full) begin // @[Reg.scala 17:18]
      victim_1Hidx_r <= _victim_1Hidx_T_2; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  victim_1Hidx = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  victim_1Hidx_r = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module L1TagAccess(
  input         clock,
  input         reset,
  input         io_r_req_valid,
  input  [4:0]  io_r_req_bits_setIdx,
  input  [21:0] io_tagFromCore_st1,
  input         io_coreReqReady,
  input         io_w_req_valid,
  input  [4:0]  io_w_req_bits_setIdx,
  input  [21:0] io_w_req_bits_data_0,
  input  [21:0] io_w_req_bits_data_1,
  output [1:0]  io_waymaskReplacement,
  output [1:0]  io_waymaskHit_st1,
  output        io_hit_st1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  wire  tagBodyAccess_clock; // @[L1CacheSubModules.scala 38:29]
  wire  tagBodyAccess_reset; // @[L1CacheSubModules.scala 38:29]
  wire  tagBodyAccess_io_r_req_valid; // @[L1CacheSubModules.scala 38:29]
  wire [4:0] tagBodyAccess_io_r_req_bits_setIdx; // @[L1CacheSubModules.scala 38:29]
  wire [21:0] tagBodyAccess_io_r_resp_data_0; // @[L1CacheSubModules.scala 38:29]
  wire [21:0] tagBodyAccess_io_r_resp_data_1; // @[L1CacheSubModules.scala 38:29]
  wire  tagBodyAccess_io_w_req_valid; // @[L1CacheSubModules.scala 38:29]
  wire [4:0] tagBodyAccess_io_w_req_bits_setIdx; // @[L1CacheSubModules.scala 38:29]
  wire [21:0] tagBodyAccess_io_w_req_bits_data_0; // @[L1CacheSubModules.scala 38:29]
  wire [21:0] tagBodyAccess_io_w_req_bits_data_1; // @[L1CacheSubModules.scala 38:29]
  wire [1:0] tagBodyAccess_io_w_req_bits_waymask; // @[L1CacheSubModules.scala 38:29]
  wire  iTagChecker_clock; // @[L1CacheSubModules.scala 53:27]
  wire  iTagChecker_reset; // @[L1CacheSubModules.scala 53:27]
  wire [21:0] iTagChecker_io_tag_of_set_0; // @[L1CacheSubModules.scala 53:27]
  wire [21:0] iTagChecker_io_tag_of_set_1; // @[L1CacheSubModules.scala 53:27]
  wire [21:0] iTagChecker_io_tag_from_pipe; // @[L1CacheSubModules.scala 53:27]
  wire  iTagChecker_io_way_valid_0; // @[L1CacheSubModules.scala 53:27]
  wire  iTagChecker_io_way_valid_1; // @[L1CacheSubModules.scala 53:27]
  wire [1:0] iTagChecker_io_waymask; // @[L1CacheSubModules.scala 53:27]
  wire  iTagChecker_io_cache_hit; // @[L1CacheSubModules.scala 53:27]
  wire  Replacement_clock; // @[L1CacheSubModules.scala 61:27]
  wire  Replacement_reset; // @[L1CacheSubModules.scala 61:27]
  wire [1:0] Replacement_io_validbits_of_set; // @[L1CacheSubModules.scala 61:27]
  wire [1:0] Replacement_io_waymask; // @[L1CacheSubModules.scala 61:27]
  wire  Replacement_io_Set_is_full; // @[L1CacheSubModules.scala 61:27]
  reg  way_valid_0_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_0_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_1_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_1_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_2_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_2_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_3_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_3_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_4_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_4_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_5_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_5_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_6_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_6_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_7_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_7_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_8_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_8_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_9_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_9_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_10_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_10_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_11_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_11_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_12_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_12_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_13_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_13_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_14_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_14_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_15_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_15_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_16_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_16_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_17_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_17_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_18_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_18_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_19_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_19_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_20_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_20_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_21_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_21_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_22_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_22_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_23_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_23_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_24_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_24_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_25_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_25_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_26_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_26_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_27_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_27_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_28_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_28_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_29_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_29_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_30_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_30_1; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_31_0; // @[L1CacheSubModules.scala 49:26]
  reg  way_valid_31_1; // @[L1CacheSubModules.scala 49:26]
  reg [4:0] iTagChecker_io_way_valid_r; // @[Reg.scala 16:16]
  wire  _GEN_2 = 5'h1 == iTagChecker_io_way_valid_r ? way_valid_1_0 : way_valid_0_0; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_3 = 5'h2 == iTagChecker_io_way_valid_r ? way_valid_2_0 : _GEN_2; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_4 = 5'h3 == iTagChecker_io_way_valid_r ? way_valid_3_0 : _GEN_3; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_5 = 5'h4 == iTagChecker_io_way_valid_r ? way_valid_4_0 : _GEN_4; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_6 = 5'h5 == iTagChecker_io_way_valid_r ? way_valid_5_0 : _GEN_5; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_7 = 5'h6 == iTagChecker_io_way_valid_r ? way_valid_6_0 : _GEN_6; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_8 = 5'h7 == iTagChecker_io_way_valid_r ? way_valid_7_0 : _GEN_7; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_9 = 5'h8 == iTagChecker_io_way_valid_r ? way_valid_8_0 : _GEN_8; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_10 = 5'h9 == iTagChecker_io_way_valid_r ? way_valid_9_0 : _GEN_9; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_11 = 5'ha == iTagChecker_io_way_valid_r ? way_valid_10_0 : _GEN_10; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_12 = 5'hb == iTagChecker_io_way_valid_r ? way_valid_11_0 : _GEN_11; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_13 = 5'hc == iTagChecker_io_way_valid_r ? way_valid_12_0 : _GEN_12; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_14 = 5'hd == iTagChecker_io_way_valid_r ? way_valid_13_0 : _GEN_13; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_15 = 5'he == iTagChecker_io_way_valid_r ? way_valid_14_0 : _GEN_14; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_16 = 5'hf == iTagChecker_io_way_valid_r ? way_valid_15_0 : _GEN_15; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_17 = 5'h10 == iTagChecker_io_way_valid_r ? way_valid_16_0 : _GEN_16; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_18 = 5'h11 == iTagChecker_io_way_valid_r ? way_valid_17_0 : _GEN_17; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_19 = 5'h12 == iTagChecker_io_way_valid_r ? way_valid_18_0 : _GEN_18; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_20 = 5'h13 == iTagChecker_io_way_valid_r ? way_valid_19_0 : _GEN_19; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_21 = 5'h14 == iTagChecker_io_way_valid_r ? way_valid_20_0 : _GEN_20; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_22 = 5'h15 == iTagChecker_io_way_valid_r ? way_valid_21_0 : _GEN_21; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_23 = 5'h16 == iTagChecker_io_way_valid_r ? way_valid_22_0 : _GEN_22; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_24 = 5'h17 == iTagChecker_io_way_valid_r ? way_valid_23_0 : _GEN_23; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_25 = 5'h18 == iTagChecker_io_way_valid_r ? way_valid_24_0 : _GEN_24; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_26 = 5'h19 == iTagChecker_io_way_valid_r ? way_valid_25_0 : _GEN_25; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_27 = 5'h1a == iTagChecker_io_way_valid_r ? way_valid_26_0 : _GEN_26; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_28 = 5'h1b == iTagChecker_io_way_valid_r ? way_valid_27_0 : _GEN_27; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_29 = 5'h1c == iTagChecker_io_way_valid_r ? way_valid_28_0 : _GEN_28; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_30 = 5'h1d == iTagChecker_io_way_valid_r ? way_valid_29_0 : _GEN_29; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_31 = 5'h1e == iTagChecker_io_way_valid_r ? way_valid_30_0 : _GEN_30; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_34 = 5'h1 == iTagChecker_io_way_valid_r ? way_valid_1_1 : way_valid_0_1; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_35 = 5'h2 == iTagChecker_io_way_valid_r ? way_valid_2_1 : _GEN_34; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_36 = 5'h3 == iTagChecker_io_way_valid_r ? way_valid_3_1 : _GEN_35; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_37 = 5'h4 == iTagChecker_io_way_valid_r ? way_valid_4_1 : _GEN_36; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_38 = 5'h5 == iTagChecker_io_way_valid_r ? way_valid_5_1 : _GEN_37; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_39 = 5'h6 == iTagChecker_io_way_valid_r ? way_valid_6_1 : _GEN_38; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_40 = 5'h7 == iTagChecker_io_way_valid_r ? way_valid_7_1 : _GEN_39; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_41 = 5'h8 == iTagChecker_io_way_valid_r ? way_valid_8_1 : _GEN_40; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_42 = 5'h9 == iTagChecker_io_way_valid_r ? way_valid_9_1 : _GEN_41; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_43 = 5'ha == iTagChecker_io_way_valid_r ? way_valid_10_1 : _GEN_42; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_44 = 5'hb == iTagChecker_io_way_valid_r ? way_valid_11_1 : _GEN_43; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_45 = 5'hc == iTagChecker_io_way_valid_r ? way_valid_12_1 : _GEN_44; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_46 = 5'hd == iTagChecker_io_way_valid_r ? way_valid_13_1 : _GEN_45; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_47 = 5'he == iTagChecker_io_way_valid_r ? way_valid_14_1 : _GEN_46; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_48 = 5'hf == iTagChecker_io_way_valid_r ? way_valid_15_1 : _GEN_47; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_49 = 5'h10 == iTagChecker_io_way_valid_r ? way_valid_16_1 : _GEN_48; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_50 = 5'h11 == iTagChecker_io_way_valid_r ? way_valid_17_1 : _GEN_49; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_51 = 5'h12 == iTagChecker_io_way_valid_r ? way_valid_18_1 : _GEN_50; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_52 = 5'h13 == iTagChecker_io_way_valid_r ? way_valid_19_1 : _GEN_51; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_53 = 5'h14 == iTagChecker_io_way_valid_r ? way_valid_20_1 : _GEN_52; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_54 = 5'h15 == iTagChecker_io_way_valid_r ? way_valid_21_1 : _GEN_53; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_55 = 5'h16 == iTagChecker_io_way_valid_r ? way_valid_22_1 : _GEN_54; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_56 = 5'h17 == iTagChecker_io_way_valid_r ? way_valid_23_1 : _GEN_55; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_57 = 5'h18 == iTagChecker_io_way_valid_r ? way_valid_24_1 : _GEN_56; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_58 = 5'h19 == iTagChecker_io_way_valid_r ? way_valid_25_1 : _GEN_57; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_59 = 5'h1a == iTagChecker_io_way_valid_r ? way_valid_26_1 : _GEN_58; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_60 = 5'h1b == iTagChecker_io_way_valid_r ? way_valid_27_1 : _GEN_59; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_61 = 5'h1c == iTagChecker_io_way_valid_r ? way_valid_28_1 : _GEN_60; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_62 = 5'h1d == iTagChecker_io_way_valid_r ? way_valid_29_1 : _GEN_61; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_63 = 5'h1e == iTagChecker_io_way_valid_r ? way_valid_30_1 : _GEN_62; // @[L1CacheSubModules.scala 56:{28,28}]
  wire  _GEN_66 = 5'h1 == io_w_req_bits_setIdx ? way_valid_1_0 : way_valid_0_0; // @[Cat.scala 31:{58,58}]
  wire  _GEN_67 = 5'h2 == io_w_req_bits_setIdx ? way_valid_2_0 : _GEN_66; // @[Cat.scala 31:{58,58}]
  wire  _GEN_68 = 5'h3 == io_w_req_bits_setIdx ? way_valid_3_0 : _GEN_67; // @[Cat.scala 31:{58,58}]
  wire  _GEN_69 = 5'h4 == io_w_req_bits_setIdx ? way_valid_4_0 : _GEN_68; // @[Cat.scala 31:{58,58}]
  wire  _GEN_70 = 5'h5 == io_w_req_bits_setIdx ? way_valid_5_0 : _GEN_69; // @[Cat.scala 31:{58,58}]
  wire  _GEN_71 = 5'h6 == io_w_req_bits_setIdx ? way_valid_6_0 : _GEN_70; // @[Cat.scala 31:{58,58}]
  wire  _GEN_72 = 5'h7 == io_w_req_bits_setIdx ? way_valid_7_0 : _GEN_71; // @[Cat.scala 31:{58,58}]
  wire  _GEN_73 = 5'h8 == io_w_req_bits_setIdx ? way_valid_8_0 : _GEN_72; // @[Cat.scala 31:{58,58}]
  wire  _GEN_74 = 5'h9 == io_w_req_bits_setIdx ? way_valid_9_0 : _GEN_73; // @[Cat.scala 31:{58,58}]
  wire  _GEN_75 = 5'ha == io_w_req_bits_setIdx ? way_valid_10_0 : _GEN_74; // @[Cat.scala 31:{58,58}]
  wire  _GEN_76 = 5'hb == io_w_req_bits_setIdx ? way_valid_11_0 : _GEN_75; // @[Cat.scala 31:{58,58}]
  wire  _GEN_77 = 5'hc == io_w_req_bits_setIdx ? way_valid_12_0 : _GEN_76; // @[Cat.scala 31:{58,58}]
  wire  _GEN_78 = 5'hd == io_w_req_bits_setIdx ? way_valid_13_0 : _GEN_77; // @[Cat.scala 31:{58,58}]
  wire  _GEN_79 = 5'he == io_w_req_bits_setIdx ? way_valid_14_0 : _GEN_78; // @[Cat.scala 31:{58,58}]
  wire  _GEN_80 = 5'hf == io_w_req_bits_setIdx ? way_valid_15_0 : _GEN_79; // @[Cat.scala 31:{58,58}]
  wire  _GEN_81 = 5'h10 == io_w_req_bits_setIdx ? way_valid_16_0 : _GEN_80; // @[Cat.scala 31:{58,58}]
  wire  _GEN_82 = 5'h11 == io_w_req_bits_setIdx ? way_valid_17_0 : _GEN_81; // @[Cat.scala 31:{58,58}]
  wire  _GEN_83 = 5'h12 == io_w_req_bits_setIdx ? way_valid_18_0 : _GEN_82; // @[Cat.scala 31:{58,58}]
  wire  _GEN_84 = 5'h13 == io_w_req_bits_setIdx ? way_valid_19_0 : _GEN_83; // @[Cat.scala 31:{58,58}]
  wire  _GEN_85 = 5'h14 == io_w_req_bits_setIdx ? way_valid_20_0 : _GEN_84; // @[Cat.scala 31:{58,58}]
  wire  _GEN_86 = 5'h15 == io_w_req_bits_setIdx ? way_valid_21_0 : _GEN_85; // @[Cat.scala 31:{58,58}]
  wire  _GEN_87 = 5'h16 == io_w_req_bits_setIdx ? way_valid_22_0 : _GEN_86; // @[Cat.scala 31:{58,58}]
  wire  _GEN_88 = 5'h17 == io_w_req_bits_setIdx ? way_valid_23_0 : _GEN_87; // @[Cat.scala 31:{58,58}]
  wire  _GEN_89 = 5'h18 == io_w_req_bits_setIdx ? way_valid_24_0 : _GEN_88; // @[Cat.scala 31:{58,58}]
  wire  _GEN_90 = 5'h19 == io_w_req_bits_setIdx ? way_valid_25_0 : _GEN_89; // @[Cat.scala 31:{58,58}]
  wire  _GEN_91 = 5'h1a == io_w_req_bits_setIdx ? way_valid_26_0 : _GEN_90; // @[Cat.scala 31:{58,58}]
  wire  _GEN_92 = 5'h1b == io_w_req_bits_setIdx ? way_valid_27_0 : _GEN_91; // @[Cat.scala 31:{58,58}]
  wire  _GEN_93 = 5'h1c == io_w_req_bits_setIdx ? way_valid_28_0 : _GEN_92; // @[Cat.scala 31:{58,58}]
  wire  _GEN_94 = 5'h1d == io_w_req_bits_setIdx ? way_valid_29_0 : _GEN_93; // @[Cat.scala 31:{58,58}]
  wire  _GEN_95 = 5'h1e == io_w_req_bits_setIdx ? way_valid_30_0 : _GEN_94; // @[Cat.scala 31:{58,58}]
  wire  _GEN_96 = 5'h1f == io_w_req_bits_setIdx ? way_valid_31_0 : _GEN_95; // @[Cat.scala 31:{58,58}]
  wire  _GEN_98 = 5'h1 == io_w_req_bits_setIdx ? way_valid_1_1 : way_valid_0_1; // @[Cat.scala 31:{58,58}]
  wire  _GEN_99 = 5'h2 == io_w_req_bits_setIdx ? way_valid_2_1 : _GEN_98; // @[Cat.scala 31:{58,58}]
  wire  _GEN_100 = 5'h3 == io_w_req_bits_setIdx ? way_valid_3_1 : _GEN_99; // @[Cat.scala 31:{58,58}]
  wire  _GEN_101 = 5'h4 == io_w_req_bits_setIdx ? way_valid_4_1 : _GEN_100; // @[Cat.scala 31:{58,58}]
  wire  _GEN_102 = 5'h5 == io_w_req_bits_setIdx ? way_valid_5_1 : _GEN_101; // @[Cat.scala 31:{58,58}]
  wire  _GEN_103 = 5'h6 == io_w_req_bits_setIdx ? way_valid_6_1 : _GEN_102; // @[Cat.scala 31:{58,58}]
  wire  _GEN_104 = 5'h7 == io_w_req_bits_setIdx ? way_valid_7_1 : _GEN_103; // @[Cat.scala 31:{58,58}]
  wire  _GEN_105 = 5'h8 == io_w_req_bits_setIdx ? way_valid_8_1 : _GEN_104; // @[Cat.scala 31:{58,58}]
  wire  _GEN_106 = 5'h9 == io_w_req_bits_setIdx ? way_valid_9_1 : _GEN_105; // @[Cat.scala 31:{58,58}]
  wire  _GEN_107 = 5'ha == io_w_req_bits_setIdx ? way_valid_10_1 : _GEN_106; // @[Cat.scala 31:{58,58}]
  wire  _GEN_108 = 5'hb == io_w_req_bits_setIdx ? way_valid_11_1 : _GEN_107; // @[Cat.scala 31:{58,58}]
  wire  _GEN_109 = 5'hc == io_w_req_bits_setIdx ? way_valid_12_1 : _GEN_108; // @[Cat.scala 31:{58,58}]
  wire  _GEN_110 = 5'hd == io_w_req_bits_setIdx ? way_valid_13_1 : _GEN_109; // @[Cat.scala 31:{58,58}]
  wire  _GEN_111 = 5'he == io_w_req_bits_setIdx ? way_valid_14_1 : _GEN_110; // @[Cat.scala 31:{58,58}]
  wire  _GEN_112 = 5'hf == io_w_req_bits_setIdx ? way_valid_15_1 : _GEN_111; // @[Cat.scala 31:{58,58}]
  wire  _GEN_113 = 5'h10 == io_w_req_bits_setIdx ? way_valid_16_1 : _GEN_112; // @[Cat.scala 31:{58,58}]
  wire  _GEN_114 = 5'h11 == io_w_req_bits_setIdx ? way_valid_17_1 : _GEN_113; // @[Cat.scala 31:{58,58}]
  wire  _GEN_115 = 5'h12 == io_w_req_bits_setIdx ? way_valid_18_1 : _GEN_114; // @[Cat.scala 31:{58,58}]
  wire  _GEN_116 = 5'h13 == io_w_req_bits_setIdx ? way_valid_19_1 : _GEN_115; // @[Cat.scala 31:{58,58}]
  wire  _GEN_117 = 5'h14 == io_w_req_bits_setIdx ? way_valid_20_1 : _GEN_116; // @[Cat.scala 31:{58,58}]
  wire  _GEN_118 = 5'h15 == io_w_req_bits_setIdx ? way_valid_21_1 : _GEN_117; // @[Cat.scala 31:{58,58}]
  wire  _GEN_119 = 5'h16 == io_w_req_bits_setIdx ? way_valid_22_1 : _GEN_118; // @[Cat.scala 31:{58,58}]
  wire  _GEN_120 = 5'h17 == io_w_req_bits_setIdx ? way_valid_23_1 : _GEN_119; // @[Cat.scala 31:{58,58}]
  wire  _GEN_121 = 5'h18 == io_w_req_bits_setIdx ? way_valid_24_1 : _GEN_120; // @[Cat.scala 31:{58,58}]
  wire  _GEN_122 = 5'h19 == io_w_req_bits_setIdx ? way_valid_25_1 : _GEN_121; // @[Cat.scala 31:{58,58}]
  wire  _GEN_123 = 5'h1a == io_w_req_bits_setIdx ? way_valid_26_1 : _GEN_122; // @[Cat.scala 31:{58,58}]
  wire  _GEN_124 = 5'h1b == io_w_req_bits_setIdx ? way_valid_27_1 : _GEN_123; // @[Cat.scala 31:{58,58}]
  wire  _GEN_125 = 5'h1c == io_w_req_bits_setIdx ? way_valid_28_1 : _GEN_124; // @[Cat.scala 31:{58,58}]
  wire  _GEN_126 = 5'h1d == io_w_req_bits_setIdx ? way_valid_29_1 : _GEN_125; // @[Cat.scala 31:{58,58}]
  wire  _GEN_127 = 5'h1e == io_w_req_bits_setIdx ? way_valid_30_1 : _GEN_126; // @[Cat.scala 31:{58,58}]
  wire  _GEN_128 = 5'h1f == io_w_req_bits_setIdx ? way_valid_31_1 : _GEN_127; // @[Cat.scala 31:{58,58}]
  wire  _GEN_129 = 5'h0 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_0_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_130 = 5'h0 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_0_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_131 = 5'h1 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_1_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_132 = 5'h1 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_1_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_133 = 5'h2 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_2_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_134 = 5'h2 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_2_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_135 = 5'h3 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_3_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_136 = 5'h3 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_3_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_137 = 5'h4 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_4_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_138 = 5'h4 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_4_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_139 = 5'h5 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_5_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_140 = 5'h5 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_5_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_141 = 5'h6 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_6_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_142 = 5'h6 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_6_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_143 = 5'h7 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_7_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_144 = 5'h7 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_7_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_145 = 5'h8 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_8_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_146 = 5'h8 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_8_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_147 = 5'h9 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_9_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_148 = 5'h9 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_9_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_149 = 5'ha == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_10_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_150 = 5'ha == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_10_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_151 = 5'hb == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_11_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_152 = 5'hb == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_11_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_153 = 5'hc == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_12_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_154 = 5'hc == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_12_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_155 = 5'hd == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_13_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_156 = 5'hd == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_13_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_157 = 5'he == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_14_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_158 = 5'he == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_14_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_159 = 5'hf == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_15_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_160 = 5'hf == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_15_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_161 = 5'h10 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_16_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_162 = 5'h10 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_16_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_163 = 5'h11 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_17_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_164 = 5'h11 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_17_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_165 = 5'h12 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_18_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_166 = 5'h12 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_18_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_167 = 5'h13 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_19_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_168 = 5'h13 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_19_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_169 = 5'h14 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_20_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_170 = 5'h14 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_20_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_171 = 5'h15 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_21_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_172 = 5'h15 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_21_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_173 = 5'h16 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_22_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_174 = 5'h16 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_22_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_175 = 5'h17 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_23_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_176 = 5'h17 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_23_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_177 = 5'h18 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_24_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_178 = 5'h18 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_24_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_179 = 5'h19 == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_25_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_180 = 5'h19 == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_25_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_181 = 5'h1a == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_26_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_182 = 5'h1a == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_26_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_183 = 5'h1b == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_27_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_184 = 5'h1b == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_27_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_185 = 5'h1c == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_28_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_186 = 5'h1c == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_28_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_187 = 5'h1d == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_29_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_188 = 5'h1d == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_29_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_189 = 5'h1e == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_30_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_190 = 5'h1e == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_30_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_191 = 5'h1f == io_w_req_bits_setIdx & ~Replacement_io_waymask[1] | way_valid_31_0; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  wire  _GEN_192 = 5'h1f == io_w_req_bits_setIdx & Replacement_io_waymask[1] | way_valid_31_1; // @[L1CacheSubModules.scala 49:26 68:{71,71}]
  SRAMTemplate tagBodyAccess ( // @[L1CacheSubModules.scala 38:29]
    .clock(tagBodyAccess_clock),
    .reset(tagBodyAccess_reset),
    .io_r_req_valid(tagBodyAccess_io_r_req_valid),
    .io_r_req_bits_setIdx(tagBodyAccess_io_r_req_bits_setIdx),
    .io_r_resp_data_0(tagBodyAccess_io_r_resp_data_0),
    .io_r_resp_data_1(tagBodyAccess_io_r_resp_data_1),
    .io_w_req_valid(tagBodyAccess_io_w_req_valid),
    .io_w_req_bits_setIdx(tagBodyAccess_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(tagBodyAccess_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(tagBodyAccess_io_w_req_bits_data_1),
    .io_w_req_bits_waymask(tagBodyAccess_io_w_req_bits_waymask)
  );
  tagChecker iTagChecker ( // @[L1CacheSubModules.scala 53:27]
    .clock(iTagChecker_clock),
    .reset(iTagChecker_reset),
    .io_tag_of_set_0(iTagChecker_io_tag_of_set_0),
    .io_tag_of_set_1(iTagChecker_io_tag_of_set_1),
    .io_tag_from_pipe(iTagChecker_io_tag_from_pipe),
    .io_way_valid_0(iTagChecker_io_way_valid_0),
    .io_way_valid_1(iTagChecker_io_way_valid_1),
    .io_waymask(iTagChecker_io_waymask),
    .io_cache_hit(iTagChecker_io_cache_hit)
  );
  ReplacementUnit Replacement ( // @[L1CacheSubModules.scala 61:27]
    .clock(Replacement_clock),
    .reset(Replacement_reset),
    .io_validbits_of_set(Replacement_io_validbits_of_set),
    .io_waymask(Replacement_io_waymask),
    .io_Set_is_full(Replacement_io_Set_is_full)
  );
  assign io_waymaskReplacement = Replacement_io_waymask; // @[L1CacheSubModules.scala 63:25]
  assign io_waymaskHit_st1 = iTagChecker_io_waymask; // @[L1CacheSubModules.scala 57:21]
  assign io_hit_st1 = iTagChecker_io_cache_hit; // @[L1CacheSubModules.scala 58:14]
  assign tagBodyAccess_clock = clock;
  assign tagBodyAccess_reset = reset;
  assign tagBodyAccess_io_r_req_valid = io_r_req_valid; // @[L1CacheSubModules.scala 47:22]
  assign tagBodyAccess_io_r_req_bits_setIdx = io_r_req_bits_setIdx; // @[L1CacheSubModules.scala 47:22]
  assign tagBodyAccess_io_w_req_valid = io_w_req_valid; // @[L1CacheSubModules.scala 64:32]
  assign tagBodyAccess_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[SRAMTemplate.scala 42:17]
  assign tagBodyAccess_io_w_req_bits_data_0 = io_w_req_bits_data_0; // @[SRAMTemplate.scala 53:15]
  assign tagBodyAccess_io_w_req_bits_data_1 = io_w_req_bits_data_1; // @[SRAMTemplate.scala 53:15]
  assign tagBodyAccess_io_w_req_bits_waymask = Replacement_io_waymask; // @[SRAMTemplate.scala 54:24]
  assign iTagChecker_clock = clock;
  assign iTagChecker_reset = reset;
  assign iTagChecker_io_tag_of_set_0 = tagBodyAccess_io_r_resp_data_0; // @[L1CacheSubModules.scala 54:29]
  assign iTagChecker_io_tag_of_set_1 = tagBodyAccess_io_r_resp_data_1; // @[L1CacheSubModules.scala 54:29]
  assign iTagChecker_io_tag_from_pipe = io_tagFromCore_st1; // @[L1CacheSubModules.scala 55:32]
  assign iTagChecker_io_way_valid_0 = 5'h1f == iTagChecker_io_way_valid_r ? way_valid_31_0 : _GEN_31; // @[L1CacheSubModules.scala 56:{28,28}]
  assign iTagChecker_io_way_valid_1 = 5'h1f == iTagChecker_io_way_valid_r ? way_valid_31_1 : _GEN_63; // @[L1CacheSubModules.scala 56:{28,28}]
  assign Replacement_clock = clock;
  assign Replacement_reset = reset;
  assign Replacement_io_validbits_of_set = {_GEN_96,_GEN_128}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_0_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_0_0 <= _GEN_129;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_0_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_0_1 <= _GEN_130;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_1_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_1_0 <= _GEN_131;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_1_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_1_1 <= _GEN_132;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_2_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_2_0 <= _GEN_133;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_2_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_2_1 <= _GEN_134;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_3_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_3_0 <= _GEN_135;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_3_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_3_1 <= _GEN_136;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_4_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_4_0 <= _GEN_137;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_4_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_4_1 <= _GEN_138;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_5_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_5_0 <= _GEN_139;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_5_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_5_1 <= _GEN_140;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_6_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_6_0 <= _GEN_141;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_6_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_6_1 <= _GEN_142;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_7_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_7_0 <= _GEN_143;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_7_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_7_1 <= _GEN_144;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_8_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_8_0 <= _GEN_145;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_8_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_8_1 <= _GEN_146;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_9_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_9_0 <= _GEN_147;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_9_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_9_1 <= _GEN_148;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_10_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_10_0 <= _GEN_149;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_10_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_10_1 <= _GEN_150;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_11_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_11_0 <= _GEN_151;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_11_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_11_1 <= _GEN_152;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_12_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_12_0 <= _GEN_153;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_12_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_12_1 <= _GEN_154;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_13_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_13_0 <= _GEN_155;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_13_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_13_1 <= _GEN_156;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_14_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_14_0 <= _GEN_157;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_14_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_14_1 <= _GEN_158;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_15_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_15_0 <= _GEN_159;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_15_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_15_1 <= _GEN_160;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_16_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_16_0 <= _GEN_161;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_16_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_16_1 <= _GEN_162;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_17_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_17_0 <= _GEN_163;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_17_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_17_1 <= _GEN_164;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_18_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_18_0 <= _GEN_165;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_18_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_18_1 <= _GEN_166;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_19_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_19_0 <= _GEN_167;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_19_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_19_1 <= _GEN_168;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_20_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_20_0 <= _GEN_169;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_20_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_20_1 <= _GEN_170;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_21_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_21_0 <= _GEN_171;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_21_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_21_1 <= _GEN_172;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_22_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_22_0 <= _GEN_173;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_22_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_22_1 <= _GEN_174;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_23_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_23_0 <= _GEN_175;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_23_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_23_1 <= _GEN_176;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_24_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_24_0 <= _GEN_177;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_24_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_24_1 <= _GEN_178;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_25_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_25_0 <= _GEN_179;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_25_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_25_1 <= _GEN_180;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_26_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_26_0 <= _GEN_181;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_26_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_26_1 <= _GEN_182;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_27_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_27_0 <= _GEN_183;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_27_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_27_1 <= _GEN_184;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_28_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_28_0 <= _GEN_185;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_28_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_28_1 <= _GEN_186;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_29_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_29_0 <= _GEN_187;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_29_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_29_1 <= _GEN_188;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_30_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_30_0 <= _GEN_189;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_30_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_30_1 <= _GEN_190;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_31_0 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_31_0 <= _GEN_191;
    end
    if (reset) begin // @[L1CacheSubModules.scala 49:26]
      way_valid_31_1 <= 1'h0; // @[L1CacheSubModules.scala 49:26]
    end else if (io_w_req_valid & ~Replacement_io_Set_is_full) begin // @[L1CacheSubModules.scala 67:54]
      way_valid_31_1 <= _GEN_192;
    end
    if (io_coreReqReady) begin // @[Reg.scala 17:18]
      iTagChecker_io_way_valid_r <= io_r_req_bits_setIdx; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  way_valid_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  way_valid_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  way_valid_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  way_valid_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  way_valid_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  way_valid_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  way_valid_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  way_valid_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  way_valid_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  way_valid_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  way_valid_5_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  way_valid_5_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  way_valid_6_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  way_valid_6_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  way_valid_7_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  way_valid_7_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  way_valid_8_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  way_valid_8_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  way_valid_9_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  way_valid_9_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_valid_10_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  way_valid_10_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  way_valid_11_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_valid_11_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_valid_12_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_valid_12_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_valid_13_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_valid_13_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_valid_14_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_valid_14_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_valid_15_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_valid_15_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_valid_16_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_valid_16_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_valid_17_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_valid_17_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_valid_18_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_valid_18_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_valid_19_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_valid_19_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_valid_20_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_valid_20_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_valid_21_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_valid_21_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_valid_22_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_valid_22_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_valid_23_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_valid_23_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_valid_24_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_valid_24_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_valid_25_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_valid_25_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_valid_26_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_valid_26_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_valid_27_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_valid_27_1 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_valid_28_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_valid_28_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_valid_29_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_valid_29_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_valid_30_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_valid_30_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_valid_31_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_valid_31_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  iTagChecker_io_way_valid_r = _RAND_64[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_1(
  input          clock,
  input          reset,
  input          io_r_req_valid,
  input  [4:0]   io_r_req_bits_setIdx,
  output [255:0] io_r_resp_data_0,
  output [255:0] io_r_resp_data_1,
  input          io_w_req_valid,
  input  [4:0]   io_w_req_bits_setIdx,
  input  [255:0] io_w_req_bits_data_0,
  input  [255:0] io_w_req_bits_data_1,
  input  [1:0]   io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [255:0] _RAND_0;
  reg [255:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] array_0 [0:31]; // @[SRAMTemplate.scala 101:26]
  wire  array_0_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_0_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [255:0] array_0_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [255:0] array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_0_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_0_raw_rdata_en_pipe_0;
  reg [4:0] array_0_raw_rdata_addr_pipe_0;
  reg [255:0] array_1 [0:31]; // @[SRAMTemplate.scala 101:26]
  wire  array_1_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_1_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [255:0] array_1_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [255:0] array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [4:0] array_1_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_1_raw_rdata_en_pipe_0;
  reg [4:0] array_1_raw_rdata_addr_pipe_0;
  reg [63:0] bypass_wdata_lfsr; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor = bypass_wdata_lfsr[0] ^ bypass_wdata_lfsr[1] ^ bypass_wdata_lfsr[3] ^ bypass_wdata_lfsr[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_2 = {bypass_wdata_xor,bypass_wdata_lfsr[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_1; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_1 = bypass_wdata_lfsr_1[0] ^ bypass_wdata_lfsr_1[1] ^ bypass_wdata_lfsr_1[3] ^
    bypass_wdata_lfsr_1[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_6 = {bypass_wdata_xor_1,bypass_wdata_lfsr_1[63:1]}; // @[Cat.scala 31:58]
  reg  bypass_mask_need_check; // @[SRAMTemplate.scala 126:29]
  reg [4:0] bypass_mask_waddr_reg; // @[SRAMTemplate.scala 127:28]
  reg [4:0] bypass_mask_raddr_reg; // @[SRAMTemplate.scala 128:28]
  wire  _bypass_mask_bypass_T_1 = bypass_mask_need_check & bypass_mask_waddr_reg == bypass_mask_raddr_reg; // @[SRAMTemplate.scala 130:39]
  wire [1:0] _bypass_mask_bypass_T_3 = _bypass_mask_bypass_T_1 ? 2'h3 : 2'h0; // @[Bitwise.scala 74:12]
  reg [1:0] bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:76]
  wire [1:0] bypass_mask_bypass = _bypass_mask_bypass_T_3 & bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:67]
  wire [255:0] bypass_wdata_0 = {{192'd0}, bypass_wdata_lfsr}; // @[SRAMTemplate.scala 134:{58,58}]
  wire [255:0] bypass_wdata_1 = {{192'd0}, bypass_wdata_lfsr_1}; // @[SRAMTemplate.scala 134:{58,58}]
  assign array_0_raw_rdata_en = array_0_raw_rdata_en_pipe_0;
  assign array_0_raw_rdata_addr = array_0_raw_rdata_addr_pipe_0;
  assign array_0_raw_rdata_data = array_0[array_0_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_0_MPORT_data = io_w_req_bits_data_0;
  assign array_0_MPORT_addr = io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = io_w_req_bits_waymask[0];
  assign array_0_MPORT_en = io_w_req_valid;
  assign array_1_raw_rdata_en = array_1_raw_rdata_en_pipe_0;
  assign array_1_raw_rdata_addr = array_1_raw_rdata_addr_pipe_0;
  assign array_1_raw_rdata_data = array_1[array_1_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_1_MPORT_data = io_w_req_bits_data_1;
  assign array_1_MPORT_addr = io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = io_w_req_bits_waymask[1];
  assign array_1_MPORT_en = io_w_req_valid;
  assign io_r_resp_data_0 = bypass_mask_bypass[0] ? bypass_wdata_0 : array_0_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_1 = bypass_mask_bypass[1] ? bypass_wdata_1 : array_1_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_0_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_0_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_1_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_1_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr <= 64'h1;
    end else begin
      bypass_wdata_lfsr <= _bypass_wdata_lfsr_T_2;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_1 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_1 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_1 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_1 <= _bypass_wdata_lfsr_T_6;
    end
    bypass_mask_need_check <= io_r_req_valid & io_w_req_valid; // @[SRAMTemplate.scala 126:34]
    bypass_mask_waddr_reg <= io_w_req_bits_setIdx; // @[SRAMTemplate.scala 127:28]
    bypass_mask_raddr_reg <= io_r_req_bits_setIdx; // @[SRAMTemplate.scala 128:28]
    bypass_mask_bypass_REG <= io_w_req_bits_waymask; // @[SRAMTemplate.scala 130:76]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {8{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    array_0[initvar] = _RAND_0[255:0];
  _RAND_3 = {8{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    array_1[initvar] = _RAND_3[255:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_raw_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_raw_rdata_addr_pipe_0 = _RAND_2[4:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_raw_rdata_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_raw_rdata_addr_pipe_0 = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  bypass_wdata_lfsr = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  bypass_wdata_lfsr_1 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  bypass_mask_need_check = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  bypass_mask_waddr_reg = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  bypass_mask_raddr_reg = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  bypass_mask_bypass_REG = _RAND_11[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module getEntryStatus(
  input  [3:0] io_valid_list,
  output       io_full,
  output [1:0] io_next,
  output [2:0] io_used
);
  wire [1:0] _io_used_T_4 = io_valid_list[0] + io_valid_list[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _io_used_T_6 = io_valid_list[2] + io_valid_list[3]; // @[Bitwise.scala 48:55]
  wire [1:0] _io_next_T_8 = ~io_valid_list[2] ? 2'h2 : 2'h3; // @[L1CacheSubModules.scala 19:55]
  wire [1:0] _io_next_T_9 = ~io_valid_list[1] ? 2'h1 : _io_next_T_8; // @[L1CacheSubModules.scala 19:55]
  assign io_full = io_used == 3'h4; // @[L1CacheSubModules.scala 18:22]
  assign io_next = ~io_valid_list[0] ? 2'h0 : _io_next_T_9; // @[L1CacheSubModules.scala 19:55]
  assign io_used = _io_used_T_4 + _io_used_T_6; // @[Bitwise.scala 48:55]
endmodule
module MSHR(
  input         clock,
  input         reset,
  output        io_missReq_ready,
  input         io_missReq_valid,
  input  [26:0] io_missReq_bits_blockAddr,
  input  [1:0]  io_missReq_bits_targetInfo,
  output        io_missRspIn_ready,
  input         io_missRspIn_valid,
  input  [26:0] io_missRspIn_bits_blockAddr,
  output        io_missRspOut_valid,
  output [26:0] io_missRspOut_bits_blockAddr,
  input         io_miss2mem_ready,
  output        io_miss2mem_valid,
  output [26:0] io_miss2mem_bits_blockAddr,
  output [1:0]  io_miss2mem_bits_instrId
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] subentryStatus_io_valid_list; // @[ICacheMSHR.scala 76:30]
  wire  subentryStatus_io_full; // @[ICacheMSHR.scala 76:30]
  wire [1:0] subentryStatus_io_next; // @[ICacheMSHR.scala 76:30]
  wire [2:0] subentryStatus_io_used; // @[ICacheMSHR.scala 76:30]
  wire [3:0] entryStatus_io_valid_list; // @[ICacheMSHR.scala 83:27]
  wire  entryStatus_io_full; // @[ICacheMSHR.scala 83:27]
  wire [1:0] entryStatus_io_next; // @[ICacheMSHR.scala 83:27]
  wire [2:0] entryStatus_io_used; // @[ICacheMSHR.scala 83:27]
  wire [3:0] hasSendStatus_io_valid_list; // @[ICacheMSHR.scala 148:29]
  wire  hasSendStatus_io_full; // @[ICacheMSHR.scala 148:29]
  wire [1:0] hasSendStatus_io_next; // @[ICacheMSHR.scala 148:29]
  wire [2:0] hasSendStatus_io_used; // @[ICacheMSHR.scala 148:29]
  reg [26:0] blockAddr_Access_0; // @[ICacheMSHR.scala 54:33]
  reg [26:0] blockAddr_Access_1; // @[ICacheMSHR.scala 54:33]
  reg [26:0] blockAddr_Access_2; // @[ICacheMSHR.scala 54:33]
  reg [26:0] blockAddr_Access_3; // @[ICacheMSHR.scala 54:33]
  reg [1:0] targetInfo_Accesss_0_0; // @[ICacheMSHR.scala 55:35]
  reg [1:0] targetInfo_Accesss_1_0; // @[ICacheMSHR.scala 55:35]
  reg [1:0] targetInfo_Accesss_2_0; // @[ICacheMSHR.scala 55:35]
  reg [1:0] targetInfo_Accesss_3_0; // @[ICacheMSHR.scala 55:35]
  reg  subentry_valid_0_0; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_0_1; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_0_2; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_0_3; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_1_0; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_1_1; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_1_2; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_1_3; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_2_0; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_2_1; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_2_2; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_2_3; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_3_0; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_3_1; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_3_2; // @[ICacheMSHR.scala 74:31]
  reg  subentry_valid_3_3; // @[ICacheMSHR.scala 74:31]
  wire  _entryMatchMissRsp_T = blockAddr_Access_0 == io_missRspIn_bits_blockAddr; // @[ICacheMSHR.scala 86:58]
  wire  _entryMatchMissRsp_T_1 = blockAddr_Access_1 == io_missRspIn_bits_blockAddr; // @[ICacheMSHR.scala 86:58]
  wire  _entryMatchMissRsp_T_2 = blockAddr_Access_2 == io_missRspIn_bits_blockAddr; // @[ICacheMSHR.scala 86:58]
  wire  _entryMatchMissRsp_T_3 = blockAddr_Access_3 == io_missRspIn_bits_blockAddr; // @[ICacheMSHR.scala 86:58]
  wire [3:0] _entryMatchMissRsp_T_4 = {_entryMatchMissRsp_T,_entryMatchMissRsp_T_1,_entryMatchMissRsp_T_2,
    _entryMatchMissRsp_T_3}; // @[Cat.scala 31:58]
  wire [3:0] _entryMatchMissRsp_T_13 = {_entryMatchMissRsp_T_4[0],_entryMatchMissRsp_T_4[1],_entryMatchMissRsp_T_4[2],
    _entryMatchMissRsp_T_4[3]}; // @[Cat.scala 31:58]
  wire [3:0] _entry_valid_T = {subentry_valid_0_0,subentry_valid_0_1,subentry_valid_0_2,subentry_valid_0_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_1 = |_entry_valid_T; // @[ICacheMSHR.scala 82:59]
  wire [3:0] _entry_valid_T_2 = {subentry_valid_1_0,subentry_valid_1_1,subentry_valid_1_2,subentry_valid_1_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_3 = |_entry_valid_T_2; // @[ICacheMSHR.scala 82:59]
  wire [3:0] _entry_valid_T_4 = {subentry_valid_2_0,subentry_valid_2_1,subentry_valid_2_2,subentry_valid_2_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_5 = |_entry_valid_T_4; // @[ICacheMSHR.scala 82:59]
  wire [3:0] _entry_valid_T_6 = {subentry_valid_3_0,subentry_valid_3_1,subentry_valid_3_2,subentry_valid_3_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_7 = |_entry_valid_T_6; // @[ICacheMSHR.scala 82:59]
  wire [3:0] _entry_valid_T_8 = {_entry_valid_T_1,_entry_valid_T_3,_entry_valid_T_5,_entry_valid_T_7}; // @[Cat.scala 31:58]
  wire [1:0] _entry_valid_T_12 = {_entry_valid_T_8[0],_entry_valid_T_8[1]}; // @[Cat.scala 31:58]
  wire [1:0] _entry_valid_T_16 = {_entry_valid_T_8[2],_entry_valid_T_8[3]}; // @[Cat.scala 31:58]
  wire [3:0] entry_valid = {_entry_valid_T_8[0],_entry_valid_T_8[1],_entry_valid_T_8[2],_entry_valid_T_8[3]}; // @[Cat.scala 31:58]
  wire [3:0] entryMatchMissRsp = _entryMatchMissRsp_T_13 & entry_valid; // @[ICacheMSHR.scala 86:92]
  wire [1:0] subentry_selected_hi = entryMatchMissRsp[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] subentry_selected_lo = entryMatchMissRsp[1:0]; // @[OneHot.scala 31:18]
  wire  _subentry_selected_T = |subentry_selected_hi; // @[OneHot.scala 32:14]
  wire [1:0] _subentry_selected_T_1 = subentry_selected_hi | subentry_selected_lo; // @[OneHot.scala 32:28]
  wire [1:0] _subentry_selected_T_3 = {_subentry_selected_T,_subentry_selected_T_1[1]}; // @[Cat.scala 31:58]
  wire  _GEN_1 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_2 : subentry_valid_0_2; // @[Cat.scala 31:{58,58}]
  wire  _GEN_2 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_2 : _GEN_1; // @[Cat.scala 31:{58,58}]
  wire  _GEN_3 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_2 : _GEN_2; // @[Cat.scala 31:{58,58}]
  wire  _GEN_5 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_3 : subentry_valid_0_3; // @[Cat.scala 31:{58,58}]
  wire  _GEN_6 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_3 : _GEN_5; // @[Cat.scala 31:{58,58}]
  wire  _GEN_7 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_3 : _GEN_6; // @[Cat.scala 31:{58,58}]
  wire  _GEN_9 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_0 : subentry_valid_0_0; // @[Cat.scala 31:{58,58}]
  wire  _GEN_10 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_0 : _GEN_9; // @[Cat.scala 31:{58,58}]
  wire  _GEN_11 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_0 : _GEN_10; // @[Cat.scala 31:{58,58}]
  wire  _GEN_13 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_1 : subentry_valid_0_1; // @[Cat.scala 31:{58,58}]
  wire  _GEN_14 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_1 : _GEN_13; // @[Cat.scala 31:{58,58}]
  wire  _GEN_15 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_1 : _GEN_14; // @[Cat.scala 31:{58,58}]
  wire [3:0] _subentryStatus_io_valid_list_T = {_GEN_11,_GEN_15,_GEN_3,_GEN_7}; // @[Cat.scala 31:58]
  wire [1:0] _subentryStatus_io_valid_list_T_4 = {_subentryStatus_io_valid_list_T[0],_subentryStatus_io_valid_list_T[1]}
    ; // @[Cat.scala 31:58]
  wire [1:0] _subentryStatus_io_valid_list_T_8 = {_subentryStatus_io_valid_list_T[2],_subentryStatus_io_valid_list_T[3]}
    ; // @[Cat.scala 31:58]
  wire [1:0] _subentry_next2cancel_T_4 = _GEN_3 ? 2'h2 : 2'h3; // @[ICacheMSHR.scala 79:55]
  wire [1:0] _subentry_next2cancel_T_5 = _GEN_15 ? 2'h1 : _subentry_next2cancel_T_4; // @[ICacheMSHR.scala 79:55]
  wire [1:0] subentry_next2cancel = _GEN_11 ? 2'h0 : _subentry_next2cancel_T_5; // @[ICacheMSHR.scala 79:55]
  wire [1:0] _T_4 = entryMatchMissRsp[0] + entryMatchMissRsp[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _T_6 = entryMatchMissRsp[2] + entryMatchMissRsp[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _T_8 = _T_4 + _T_6; // @[Bitwise.scala 48:55]
  wire  _T_12 = ~reset; // @[ICacheMSHR.scala 87:9]
  wire  _entryMatchMissReq_T = blockAddr_Access_0 == io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 88:58]
  wire  _entryMatchMissReq_T_1 = blockAddr_Access_1 == io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 88:58]
  wire  _entryMatchMissReq_T_2 = blockAddr_Access_2 == io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 88:58]
  wire  _entryMatchMissReq_T_3 = blockAddr_Access_3 == io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 88:58]
  wire [3:0] _entryMatchMissReq_T_4 = {_entryMatchMissReq_T,_entryMatchMissReq_T_1,_entryMatchMissReq_T_2,
    _entryMatchMissReq_T_3}; // @[Cat.scala 31:58]
  wire [3:0] _entryMatchMissReq_T_13 = {_entryMatchMissReq_T_4[0],_entryMatchMissReq_T_4[1],_entryMatchMissReq_T_4[2],
    _entryMatchMissReq_T_4[3]}; // @[Cat.scala 31:58]
  wire [3:0] entryMatchMissReq = _entryMatchMissReq_T_13 & entry_valid; // @[ICacheMSHR.scala 88:90]
  wire [1:0] _T_18 = entryMatchMissReq[0] + entryMatchMissReq[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _T_20 = entryMatchMissReq[2] + entryMatchMissReq[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _T_22 = _T_18 + _T_20; // @[Bitwise.scala 48:55]
  wire  secondary_miss = |entryMatchMissReq; // @[ICacheMSHR.scala 91:42]
  wire  primary_miss = ~secondary_miss; // @[ICacheMSHR.scala 92:22]
  reg  missRsqBusy; // @[ICacheMSHR.scala 95:28]
  wire  _io_missReq_ready_T_1 = subentryStatus_io_full & secondary_miss; // @[ICacheMSHR.scala 98:29]
  wire  _io_missReq_ready_T_2 = entryStatus_io_full & primary_miss | _io_missReq_ready_T_1; // @[ICacheMSHR.scala 97:63]
  wire  _ReqConflictWithRsp_T = io_missRspIn_ready & io_missRspIn_valid; // @[Decoupled.scala 50:35]
  wire  _ReqConflictWithRsp_T_4 = missRsqBusy & io_missRspOut_bits_blockAddr == io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 167:20]
  wire  _ReqConflictWithRsp_T_5 = _ReqConflictWithRsp_T & io_missRspIn_bits_blockAddr == io_missReq_bits_blockAddr |
    _ReqConflictWithRsp_T_4; // @[ICacheMSHR.scala 166:89]
  wire  ReqConflictWithRsp = io_missReq_valid & _ReqConflictWithRsp_T_5; // @[ICacheMSHR.scala 165:42]
  wire  _io_missReq_ready_T_3 = _io_missReq_ready_T_2 | ReqConflictWithRsp; // @[ICacheMSHR.scala 98:48]
  wire [1:0] tAEntryIdx_hi = entryMatchMissReq[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] tAEntryIdx_lo = entryMatchMissReq[1:0]; // @[OneHot.scala 31:18]
  wire  _tAEntryIdx_T = |tAEntryIdx_hi; // @[OneHot.scala 32:14]
  wire [1:0] _tAEntryIdx_T_1 = tAEntryIdx_hi | tAEntryIdx_lo; // @[OneHot.scala 32:28]
  wire [1:0] _tAEntryIdx_T_3 = {_tAEntryIdx_T,_tAEntryIdx_T_1[1]}; // @[Cat.scala 31:58]
  wire [1:0] tAEntryIdx = secondary_miss ? _tAEntryIdx_T_3 : entryStatus_io_next; // @[ICacheMSHR.scala 100:23]
  wire [1:0] tASubEntryIdx = secondary_miss ? subentryStatus_io_next : 2'h0; // @[ICacheMSHR.scala 101:26]
  wire  _T_28 = io_missReq_ready & io_missReq_valid; // @[Decoupled.scala 50:35]
  wire  _T_43 = subentryStatus_io_used == 3'h1; // @[ICacheMSHR.scala 112:52]
  wire  _GEN_48 = missRsqBusy & subentryStatus_io_used == 3'h1 ? 1'h0 : missRsqBusy; // @[ICacheMSHR.scala 112:83 113:17 95:28]
  wire  _GEN_49 = _ReqConflictWithRsp_T & subentryStatus_io_used != 3'h1 | _GEN_48; // @[ICacheMSHR.scala 110:88 111:17]
  wire  _GEN_196 = 2'h0 == _subentry_selected_T_3; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_197 = 2'h1 == subentry_next2cancel; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_199 = 2'h2 == subentry_next2cancel; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_201 = 2'h3 == subentry_next2cancel; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_202 = 2'h1 == _subentry_selected_T_3; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_203 = 2'h0 == subentry_next2cancel; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_210 = 2'h2 == _subentry_selected_T_3; // @[ICacheMSHR.scala 119:{33,33}]
  wire  _GEN_218 = 2'h3 == _subentry_selected_T_3; // @[ICacheMSHR.scala 119:{33,33}]
  wire [26:0] _GEN_67 = 2'h1 == _subentry_selected_T_3 ? blockAddr_Access_1 : blockAddr_Access_0; // @[ICacheMSHR.scala 120:{32,32}]
  wire [26:0] _GEN_68 = 2'h2 == _subentry_selected_T_3 ? blockAddr_Access_2 : _GEN_67; // @[ICacheMSHR.scala 120:{32,32}]
  wire  _T_47 = 2'h0 == entryStatus_io_next; // @[ICacheMSHR.scala 126:26]
  wire  _T_56 = 2'h0 == subentryStatus_io_next; // @[ICacheMSHR.scala 130:26]
  wire  _T_57 = 2'h0 == _tAEntryIdx_T_3 & _T_56; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_70 = _T_57 & secondary_miss | subentry_valid_0_0; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _GEN_71 = _T_47 & primary_miss | _GEN_70; // @[ICacheMSHR.scala 127:49 128:43]
  wire  _T_65 = io_missRspOut_valid & _GEN_196; // @[ICacheMSHR.scala 133:39]
  wire  _T_67 = _T_65 & _GEN_203; // @[ICacheMSHR.scala 134:52]
  wire  _T_78 = 2'h1 == subentryStatus_io_next; // @[ICacheMSHR.scala 130:26]
  wire  _T_79 = 2'h0 == _tAEntryIdx_T_3 & _T_78; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_74 = _T_79 & secondary_miss | subentry_valid_0_1; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_89 = _T_65 & _GEN_197; // @[ICacheMSHR.scala 134:52]
  wire  _T_100 = 2'h2 == subentryStatus_io_next; // @[ICacheMSHR.scala 130:26]
  wire  _T_101 = 2'h0 == _tAEntryIdx_T_3 & _T_100; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_78 = _T_101 & secondary_miss | subentry_valid_0_2; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_111 = _T_65 & _GEN_199; // @[ICacheMSHR.scala 134:52]
  wire  _T_122 = 2'h3 == subentryStatus_io_next; // @[ICacheMSHR.scala 130:26]
  wire  _T_123 = 2'h0 == _tAEntryIdx_T_3 & _T_122; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_82 = _T_123 & secondary_miss | subentry_valid_0_3; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_133 = _T_65 & _GEN_201; // @[ICacheMSHR.scala 134:52]
  wire  _T_135 = 2'h1 == entryStatus_io_next; // @[ICacheMSHR.scala 126:26]
  wire  _T_145 = 2'h1 == _tAEntryIdx_T_3 & _T_56; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_86 = _T_145 & secondary_miss | subentry_valid_1_0; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _GEN_87 = _T_135 & primary_miss | _GEN_86; // @[ICacheMSHR.scala 127:49 128:43]
  wire  _T_153 = io_missRspOut_valid & _GEN_202; // @[ICacheMSHR.scala 133:39]
  wire  _T_155 = _T_153 & _GEN_203; // @[ICacheMSHR.scala 134:52]
  wire  _T_167 = 2'h1 == _tAEntryIdx_T_3 & _T_78; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_90 = _T_167 & secondary_miss | subentry_valid_1_1; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_177 = _T_153 & _GEN_197; // @[ICacheMSHR.scala 134:52]
  wire  _T_189 = 2'h1 == _tAEntryIdx_T_3 & _T_100; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_94 = _T_189 & secondary_miss | subentry_valid_1_2; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_199 = _T_153 & _GEN_199; // @[ICacheMSHR.scala 134:52]
  wire  _T_211 = 2'h1 == _tAEntryIdx_T_3 & _T_122; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_98 = _T_211 & secondary_miss | subentry_valid_1_3; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_221 = _T_153 & _GEN_201; // @[ICacheMSHR.scala 134:52]
  wire  _T_223 = 2'h2 == entryStatus_io_next; // @[ICacheMSHR.scala 126:26]
  wire  _T_233 = 2'h2 == _tAEntryIdx_T_3 & _T_56; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_102 = _T_233 & secondary_miss | subentry_valid_2_0; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _GEN_103 = _T_223 & primary_miss | _GEN_102; // @[ICacheMSHR.scala 127:49 128:43]
  wire  _T_241 = io_missRspOut_valid & _GEN_210; // @[ICacheMSHR.scala 133:39]
  wire  _T_243 = _T_241 & _GEN_203; // @[ICacheMSHR.scala 134:52]
  wire  _T_255 = 2'h2 == _tAEntryIdx_T_3 & _T_78; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_106 = _T_255 & secondary_miss | subentry_valid_2_1; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_265 = _T_241 & _GEN_197; // @[ICacheMSHR.scala 134:52]
  wire  _T_277 = 2'h2 == _tAEntryIdx_T_3 & _T_100; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_110 = _T_277 & secondary_miss | subentry_valid_2_2; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_287 = _T_241 & _GEN_199; // @[ICacheMSHR.scala 134:52]
  wire  _T_299 = 2'h2 == _tAEntryIdx_T_3 & _T_122; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_114 = _T_299 & secondary_miss | subentry_valid_2_3; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_309 = _T_241 & _GEN_201; // @[ICacheMSHR.scala 134:52]
  wire  _T_311 = 2'h3 == entryStatus_io_next; // @[ICacheMSHR.scala 126:26]
  wire  _T_321 = 2'h3 == _tAEntryIdx_T_3 & _T_56; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_118 = _T_321 & secondary_miss | subentry_valid_3_0; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _GEN_119 = _T_311 & primary_miss | _GEN_118; // @[ICacheMSHR.scala 127:49 128:43]
  wire  _T_329 = io_missRspOut_valid & _GEN_218; // @[ICacheMSHR.scala 133:39]
  wire  _T_331 = _T_329 & _GEN_203; // @[ICacheMSHR.scala 134:52]
  wire  _T_343 = 2'h3 == _tAEntryIdx_T_3 & _T_78; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_122 = _T_343 & secondary_miss | subentry_valid_3_1; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_353 = _T_329 & _GEN_197; // @[ICacheMSHR.scala 134:52]
  wire  _T_365 = 2'h3 == _tAEntryIdx_T_3 & _T_100; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_126 = _T_365 & secondary_miss | subentry_valid_3_2; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_375 = _T_329 & _GEN_199; // @[ICacheMSHR.scala 134:52]
  wire  _T_387 = 2'h3 == _tAEntryIdx_T_3 & _T_122; // @[ICacheMSHR.scala 129:63]
  wire  _GEN_130 = _T_387 & secondary_miss | subentry_valid_3_3; // @[ICacheMSHR.scala 130:70 131:43 74:31]
  wire  _T_397 = _T_329 & _GEN_201; // @[ICacheMSHR.scala 134:52]
  reg  has_send2mem_0; // @[ICacheMSHR.scala 147:29]
  reg  has_send2mem_1; // @[ICacheMSHR.scala 147:29]
  reg  has_send2mem_2; // @[ICacheMSHR.scala 147:29]
  reg  has_send2mem_3; // @[ICacheMSHR.scala 147:29]
  wire [3:0] _hasSendStatus_io_valid_list_T = {has_send2mem_0,has_send2mem_1,has_send2mem_2,has_send2mem_3}; // @[Cat.scala 31:58]
  wire [1:0] _hasSendStatus_io_valid_list_T_4 = {_hasSendStatus_io_valid_list_T[0],_hasSendStatus_io_valid_list_T[1]}; // @[Cat.scala 31:58]
  wire [1:0] _hasSendStatus_io_valid_list_T_8 = {_hasSendStatus_io_valid_list_T[2],_hasSendStatus_io_valid_list_T[3]}; // @[Cat.scala 31:58]
  wire  _GEN_143 = 2'h1 == hasSendStatus_io_next ? has_send2mem_1 : has_send2mem_0; // @[ICacheMSHR.scala 150:{24,24}]
  wire  _GEN_144 = 2'h2 == hasSendStatus_io_next ? has_send2mem_2 : _GEN_143; // @[ICacheMSHR.scala 150:{24,24}]
  wire  _GEN_145 = 2'h3 == hasSendStatus_io_next ? has_send2mem_3 : _GEN_144; // @[ICacheMSHR.scala 150:{24,24}]
  wire [3:0] _io_miss2mem_valid_T_1 = entry_valid >> hasSendStatus_io_next; // @[ICacheMSHR.scala 150:75]
  wire  miss2mem_fire = io_miss2mem_valid & io_miss2mem_ready; // @[ICacheMSHR.scala 151:41]
  wire  _GEN_146 = (missRsqBusy | _ReqConflictWithRsp_T) & io_missRspOut_valid & _T_43 & _GEN_196 ? 1'h0 :
    has_send2mem_0; // @[ICacheMSHR.scala 156:146 157:25 147:29]
  wire  _GEN_147 = miss2mem_fire & 2'h0 == hasSendStatus_io_next | _GEN_146; // @[ICacheMSHR.scala 154:57 155:25]
  wire  _GEN_148 = (missRsqBusy | _ReqConflictWithRsp_T) & io_missRspOut_valid & _T_43 & _GEN_202 ? 1'h0 :
    has_send2mem_1; // @[ICacheMSHR.scala 156:146 157:25 147:29]
  wire  _GEN_149 = miss2mem_fire & 2'h1 == hasSendStatus_io_next | _GEN_148; // @[ICacheMSHR.scala 154:57 155:25]
  wire  _GEN_150 = (missRsqBusy | _ReqConflictWithRsp_T) & io_missRspOut_valid & _T_43 & _GEN_210 ? 1'h0 :
    has_send2mem_2; // @[ICacheMSHR.scala 156:146 157:25 147:29]
  wire  _GEN_151 = miss2mem_fire & 2'h2 == hasSendStatus_io_next | _GEN_150; // @[ICacheMSHR.scala 154:57 155:25]
  wire  _GEN_152 = (missRsqBusy | _ReqConflictWithRsp_T) & io_missRspOut_valid & _T_43 & _GEN_218 ? 1'h0 :
    has_send2mem_3; // @[ICacheMSHR.scala 156:146 157:25 147:29]
  wire  _GEN_153 = miss2mem_fire & 2'h3 == hasSendStatus_io_next | _GEN_152; // @[ICacheMSHR.scala 154:57 155:25]
  wire [2:0] _GEN_226 = {{1'd0}, hasSendStatus_io_next}; // @[ICacheMSHR.scala 154:31]
  wire [2:0] _GEN_227 = {{1'd0}, _subentry_selected_T_3}; // @[ICacheMSHR.scala 156:114]
  wire  _GEN_154 = (missRsqBusy | _ReqConflictWithRsp_T) & io_missRspOut_valid & _T_43 & 3'h4 == _GEN_227 ? 1'h0 :
    _GEN_147; // @[ICacheMSHR.scala 156:146 157:25]
  wire  _GEN_155 = miss2mem_fire & 3'h4 == _GEN_226 | _GEN_154; // @[ICacheMSHR.scala 154:57 155:25]
  wire [26:0] _GEN_157 = 2'h1 == hasSendStatus_io_next ? blockAddr_Access_1 : blockAddr_Access_0; // @[ICacheMSHR.scala 160:{30,30}]
  wire [26:0] _GEN_158 = 2'h2 == hasSendStatus_io_next ? blockAddr_Access_2 : _GEN_157; // @[ICacheMSHR.scala 160:{30,30}]
  wire [1:0] _GEN_161 = 2'h1 == hasSendStatus_io_next ? targetInfo_Accesss_1_0 : targetInfo_Accesss_0_0; // @[ICacheMSHR.scala 161:{28,28}]
  wire [1:0] _GEN_162 = 2'h2 == hasSendStatus_io_next ? targetInfo_Accesss_2_0 : _GEN_161; // @[ICacheMSHR.scala 161:{28,28}]
  getEntryStatus subentryStatus ( // @[ICacheMSHR.scala 76:30]
    .io_valid_list(subentryStatus_io_valid_list),
    .io_full(subentryStatus_io_full),
    .io_next(subentryStatus_io_next),
    .io_used(subentryStatus_io_used)
  );
  getEntryStatus entryStatus ( // @[ICacheMSHR.scala 83:27]
    .io_valid_list(entryStatus_io_valid_list),
    .io_full(entryStatus_io_full),
    .io_next(entryStatus_io_next),
    .io_used(entryStatus_io_used)
  );
  getEntryStatus hasSendStatus ( // @[ICacheMSHR.scala 148:29]
    .io_valid_list(hasSendStatus_io_valid_list),
    .io_full(hasSendStatus_io_full),
    .io_next(hasSendStatus_io_next),
    .io_used(hasSendStatus_io_used)
  );
  assign io_missReq_ready = ~_io_missReq_ready_T_3; // @[ICacheMSHR.scala 97:23]
  assign io_missRspIn_ready = ~missRsqBusy; // @[ICacheMSHR.scala 116:25]
  assign io_missRspOut_valid = _ReqConflictWithRsp_T | missRsqBusy; // @[ICacheMSHR.scala 117:46]
  assign io_missRspOut_bits_blockAddr = 2'h3 == _subentry_selected_T_3 ? blockAddr_Access_3 : _GEN_68; // @[ICacheMSHR.scala 120:{32,32}]
  assign io_miss2mem_valid = ~_GEN_145 & _io_miss2mem_valid_T_1[0]; // @[ICacheMSHR.scala 150:61]
  assign io_miss2mem_bits_blockAddr = 2'h3 == hasSendStatus_io_next ? blockAddr_Access_3 : _GEN_158; // @[ICacheMSHR.scala 160:{30,30}]
  assign io_miss2mem_bits_instrId = 2'h3 == hasSendStatus_io_next ? targetInfo_Accesss_3_0 : _GEN_162; // @[ICacheMSHR.scala 161:{28,28}]
  assign subentryStatus_io_valid_list = {_subentryStatus_io_valid_list_T_4,_subentryStatus_io_valid_list_T_8}; // @[Cat.scala 31:58]
  assign entryStatus_io_valid_list = {_entry_valid_T_12,_entry_valid_T_16}; // @[Cat.scala 31:58]
  assign hasSendStatus_io_valid_list = {_hasSendStatus_io_valid_list_T_4,_hasSendStatus_io_valid_list_T_8}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[ICacheMSHR.scala 54:33]
      blockAddr_Access_0 <= 27'h0; // @[ICacheMSHR.scala 54:33]
    end else if (_T_28 & primary_miss) begin // @[ICacheMSHR.scala 142:42]
      if (2'h0 == entryStatus_io_next) begin // @[ICacheMSHR.scala 143:43]
        blockAddr_Access_0 <= io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 143:43]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 54:33]
      blockAddr_Access_1 <= 27'h0; // @[ICacheMSHR.scala 54:33]
    end else if (_T_28 & primary_miss) begin // @[ICacheMSHR.scala 142:42]
      if (2'h1 == entryStatus_io_next) begin // @[ICacheMSHR.scala 143:43]
        blockAddr_Access_1 <= io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 143:43]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 54:33]
      blockAddr_Access_2 <= 27'h0; // @[ICacheMSHR.scala 54:33]
    end else if (_T_28 & primary_miss) begin // @[ICacheMSHR.scala 142:42]
      if (2'h2 == entryStatus_io_next) begin // @[ICacheMSHR.scala 143:43]
        blockAddr_Access_2 <= io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 143:43]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 54:33]
      blockAddr_Access_3 <= 27'h0; // @[ICacheMSHR.scala 54:33]
    end else if (_T_28 & primary_miss) begin // @[ICacheMSHR.scala 142:42]
      if (2'h3 == entryStatus_io_next) begin // @[ICacheMSHR.scala 143:43]
        blockAddr_Access_3 <= io_missReq_bits_blockAddr; // @[ICacheMSHR.scala 143:43]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 55:35]
      targetInfo_Accesss_0_0 <= 2'h0; // @[ICacheMSHR.scala 55:35]
    end else if (_T_28) begin // @[ICacheMSHR.scala 103:27]
      if (2'h0 == tAEntryIdx & 2'h0 == tASubEntryIdx) begin // @[ICacheMSHR.scala 104:51]
        targetInfo_Accesss_0_0 <= io_missReq_bits_targetInfo; // @[ICacheMSHR.scala 104:51]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 55:35]
      targetInfo_Accesss_1_0 <= 2'h0; // @[ICacheMSHR.scala 55:35]
    end else if (_T_28) begin // @[ICacheMSHR.scala 103:27]
      if (2'h1 == tAEntryIdx & 2'h0 == tASubEntryIdx) begin // @[ICacheMSHR.scala 104:51]
        targetInfo_Accesss_1_0 <= io_missReq_bits_targetInfo; // @[ICacheMSHR.scala 104:51]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 55:35]
      targetInfo_Accesss_2_0 <= 2'h0; // @[ICacheMSHR.scala 55:35]
    end else if (_T_28) begin // @[ICacheMSHR.scala 103:27]
      if (2'h2 == tAEntryIdx & 2'h0 == tASubEntryIdx) begin // @[ICacheMSHR.scala 104:51]
        targetInfo_Accesss_2_0 <= io_missReq_bits_targetInfo; // @[ICacheMSHR.scala 104:51]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 55:35]
      targetInfo_Accesss_3_0 <= 2'h0; // @[ICacheMSHR.scala 55:35]
    end else if (_T_28) begin // @[ICacheMSHR.scala 103:27]
      if (2'h3 == tAEntryIdx & 2'h0 == tASubEntryIdx) begin // @[ICacheMSHR.scala 104:51]
        targetInfo_Accesss_3_0 <= io_missReq_bits_targetInfo; // @[ICacheMSHR.scala 104:51]
      end
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_0_0 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_0_0 <= _GEN_71;
    end else if (_T_67) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_0_0 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_0_1 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_0_1 <= _GEN_74;
    end else if (_T_89) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_0_1 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_0_2 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_0_2 <= _GEN_78;
    end else if (_T_111) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_0_2 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_0_3 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_0_3 <= _GEN_82;
    end else if (_T_133) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_0_3 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_1_0 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_1_0 <= _GEN_87;
    end else if (_T_155) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_1_0 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_1_1 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_1_1 <= _GEN_90;
    end else if (_T_177) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_1_1 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_1_2 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_1_2 <= _GEN_94;
    end else if (_T_199) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_1_2 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_1_3 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_1_3 <= _GEN_98;
    end else if (_T_221) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_1_3 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_2_0 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_2_0 <= _GEN_103;
    end else if (_T_243) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_2_0 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_2_1 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_2_1 <= _GEN_106;
    end else if (_T_265) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_2_1 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_2_2 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_2_2 <= _GEN_110;
    end else if (_T_287) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_2_2 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_2_3 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_2_3 <= _GEN_114;
    end else if (_T_309) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_2_3 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_3_0 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_3_0 <= _GEN_119;
    end else if (_T_331) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_3_0 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_3_1 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_3_1 <= _GEN_122;
    end else if (_T_353) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_3_1 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_3_2 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_3_2 <= _GEN_126;
    end else if (_T_375) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_3_2 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 74:31]
      subentry_valid_3_3 <= 1'h0; // @[ICacheMSHR.scala 74:31]
    end else if (_T_28) begin // @[ICacheMSHR.scala 125:30]
      subentry_valid_3_3 <= _GEN_130;
    end else if (_T_397) begin // @[ICacheMSHR.scala 135:48]
      subentry_valid_3_3 <= 1'h0; // @[ICacheMSHR.scala 136:41]
    end
    if (reset) begin // @[ICacheMSHR.scala 95:28]
      missRsqBusy <= 1'h0; // @[ICacheMSHR.scala 95:28]
    end else begin
      missRsqBusy <= _GEN_49;
    end
    if (reset) begin // @[ICacheMSHR.scala 147:29]
      has_send2mem_0 <= 1'h0; // @[ICacheMSHR.scala 147:29]
    end else begin
      has_send2mem_0 <= _GEN_155;
    end
    if (reset) begin // @[ICacheMSHR.scala 147:29]
      has_send2mem_1 <= 1'h0; // @[ICacheMSHR.scala 147:29]
    end else begin
      has_send2mem_1 <= _GEN_149;
    end
    if (reset) begin // @[ICacheMSHR.scala 147:29]
      has_send2mem_2 <= 1'h0; // @[ICacheMSHR.scala 147:29]
    end else begin
      has_send2mem_2 <= _GEN_151;
    end
    if (reset) begin // @[ICacheMSHR.scala 147:29]
      has_send2mem_3 <= 1'h0; // @[ICacheMSHR.scala 147:29]
    end else begin
      has_send2mem_3 <= _GEN_153;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(_T_8 <= 3'h1)) begin
          $fatal; // @[ICacheMSHR.scala 87:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_8 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ICacheMSHR.scala:87 assert(PopCount(entryMatchMissRsp) <= 1.U)\n"); // @[ICacheMSHR.scala 87:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_12 & ~(_T_22 <= 3'h1)) begin
          $fatal; // @[ICacheMSHR.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_12 & ~(_T_22 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ICacheMSHR.scala:89 assert(PopCount(entryMatchMissReq) <= 1.U)\n"); // @[ICacheMSHR.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_12 & ~(~_ReqConflictWithRsp_T | _ReqConflictWithRsp_T & subentryStatus_io_used >= 3'h1)) begin
          $fatal; // @[ICacheMSHR.scala 108:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_12 & ~(~_ReqConflictWithRsp_T | _ReqConflictWithRsp_T & subentryStatus_io_used >= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ICacheMSHR.scala:108 assert(!io.missRspIn.fire() || (io.missRspIn.fire() && subentryStatus.io.used >= 1.U))\n"
            ); // @[ICacheMSHR.scala 108:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  blockAddr_Access_0 = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  blockAddr_Access_1 = _RAND_1[26:0];
  _RAND_2 = {1{`RANDOM}};
  blockAddr_Access_2 = _RAND_2[26:0];
  _RAND_3 = {1{`RANDOM}};
  blockAddr_Access_3 = _RAND_3[26:0];
  _RAND_4 = {1{`RANDOM}};
  targetInfo_Accesss_0_0 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  targetInfo_Accesss_1_0 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  targetInfo_Accesss_2_0 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  targetInfo_Accesss_3_0 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  subentry_valid_0_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  subentry_valid_0_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  subentry_valid_0_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  subentry_valid_0_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  subentry_valid_1_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  subentry_valid_1_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  subentry_valid_1_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  subentry_valid_1_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  subentry_valid_2_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  subentry_valid_2_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  subentry_valid_2_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  subentry_valid_2_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  subentry_valid_3_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  subentry_valid_3_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  subentry_valid_3_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  subentry_valid_3_3 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  missRsqBusy = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  has_send2mem_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  has_send2mem_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  has_send2mem_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  has_send2mem_3 = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_49(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_d_addr,
  input  [31:0] io_enq_bits_d_data_0,
  input  [31:0] io_enq_bits_d_data_1,
  input  [31:0] io_enq_bits_d_data_2,
  input  [31:0] io_enq_bits_d_data_3,
  input  [31:0] io_enq_bits_d_data_4,
  input  [31:0] io_enq_bits_d_data_5,
  input  [31:0] io_enq_bits_d_data_6,
  input  [31:0] io_enq_bits_d_data_7,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_d_addr,
  output [31:0] io_deq_bits_d_data_0,
  output [31:0] io_deq_bits_d_data_1,
  output [31:0] io_deq_bits_d_data_2,
  output [31:0] io_deq_bits_d_data_3,
  output [31:0] io_deq_bits_d_data_4,
  output [31:0] io_deq_bits_d_data_5,
  output [31:0] io_deq_bits_d_data_6,
  output [31:0] io_deq_bits_d_data_7
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_d_addr [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_addr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_addr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_addr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_addr_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_0 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_1 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_2 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_3 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_4 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_5 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_6 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_d_data_7 [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_d_data_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_d_data_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_d_data_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_d_data_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_d_data_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_d_data_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_d_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_addr_io_deq_bits_MPORT_data = ram_d_addr[ram_d_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_addr_MPORT_data = io_enq_bits_d_addr;
  assign ram_d_addr_MPORT_addr = enq_ptr_value;
  assign ram_d_addr_MPORT_mask = 1'h1;
  assign ram_d_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_0_io_deq_bits_MPORT_data = ram_d_data_0[ram_d_data_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_0_MPORT_data = io_enq_bits_d_data_0;
  assign ram_d_data_0_MPORT_addr = enq_ptr_value;
  assign ram_d_data_0_MPORT_mask = 1'h1;
  assign ram_d_data_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_1_io_deq_bits_MPORT_data = ram_d_data_1[ram_d_data_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_1_MPORT_data = io_enq_bits_d_data_1;
  assign ram_d_data_1_MPORT_addr = enq_ptr_value;
  assign ram_d_data_1_MPORT_mask = 1'h1;
  assign ram_d_data_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_2_io_deq_bits_MPORT_data = ram_d_data_2[ram_d_data_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_2_MPORT_data = io_enq_bits_d_data_2;
  assign ram_d_data_2_MPORT_addr = enq_ptr_value;
  assign ram_d_data_2_MPORT_mask = 1'h1;
  assign ram_d_data_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_3_io_deq_bits_MPORT_data = ram_d_data_3[ram_d_data_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_3_MPORT_data = io_enq_bits_d_data_3;
  assign ram_d_data_3_MPORT_addr = enq_ptr_value;
  assign ram_d_data_3_MPORT_mask = 1'h1;
  assign ram_d_data_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_4_io_deq_bits_MPORT_data = ram_d_data_4[ram_d_data_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_4_MPORT_data = io_enq_bits_d_data_4;
  assign ram_d_data_4_MPORT_addr = enq_ptr_value;
  assign ram_d_data_4_MPORT_mask = 1'h1;
  assign ram_d_data_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_5_io_deq_bits_MPORT_data = ram_d_data_5[ram_d_data_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_5_MPORT_data = io_enq_bits_d_data_5;
  assign ram_d_data_5_MPORT_addr = enq_ptr_value;
  assign ram_d_data_5_MPORT_mask = 1'h1;
  assign ram_d_data_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_6_io_deq_bits_MPORT_data = ram_d_data_6[ram_d_data_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_6_MPORT_data = io_enq_bits_d_data_6;
  assign ram_d_data_6_MPORT_addr = enq_ptr_value;
  assign ram_d_data_6_MPORT_mask = 1'h1;
  assign ram_d_data_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_d_data_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_d_data_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_d_data_7_io_deq_bits_MPORT_data = ram_d_data_7[ram_d_data_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_d_data_7_MPORT_data = io_enq_bits_d_data_7;
  assign ram_d_data_7_MPORT_addr = enq_ptr_value;
  assign ram_d_data_7_MPORT_mask = 1'h1;
  assign ram_d_data_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_d_addr = ram_d_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_0 = ram_d_data_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_1 = ram_d_data_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_2 = ram_d_data_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_3 = ram_d_data_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_4 = ram_d_data_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_5 = ram_d_data_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_6 = ram_d_data_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_d_data_7 = ram_d_data_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_d_addr_MPORT_en & ram_d_addr_MPORT_mask) begin
      ram_d_addr[ram_d_addr_MPORT_addr] <= ram_d_addr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_0_MPORT_en & ram_d_data_0_MPORT_mask) begin
      ram_d_data_0[ram_d_data_0_MPORT_addr] <= ram_d_data_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_1_MPORT_en & ram_d_data_1_MPORT_mask) begin
      ram_d_data_1[ram_d_data_1_MPORT_addr] <= ram_d_data_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_2_MPORT_en & ram_d_data_2_MPORT_mask) begin
      ram_d_data_2[ram_d_data_2_MPORT_addr] <= ram_d_data_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_3_MPORT_en & ram_d_data_3_MPORT_mask) begin
      ram_d_data_3[ram_d_data_3_MPORT_addr] <= ram_d_data_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_4_MPORT_en & ram_d_data_4_MPORT_mask) begin
      ram_d_data_4[ram_d_data_4_MPORT_addr] <= ram_d_data_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_5_MPORT_en & ram_d_data_5_MPORT_mask) begin
      ram_d_data_5[ram_d_data_5_MPORT_addr] <= ram_d_data_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_6_MPORT_en & ram_d_data_6_MPORT_mask) begin
      ram_d_data_6[ram_d_data_6_MPORT_addr] <= ram_d_data_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_d_data_7_MPORT_en & ram_d_data_7_MPORT_mask) begin
      ram_d_data_7[ram_d_data_7_MPORT_addr] <= ram_d_data_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_0[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_1[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_2[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_3[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_4[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_5[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_6[initvar] = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_d_data_7[initvar] = _RAND_8[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  enq_ptr_value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  deq_ptr_value = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  maybe_full = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstructionCache(
  input         clock,
  input         reset,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_addr,
  input  [1:0]  io_coreReq_bits_warpid,
  input         io_externalFlushPipe_valid,
  input  [1:0]  io_externalFlushPipe_bits_warpid,
  output        io_coreRsp_valid,
  output [31:0] io_coreRsp_bits_addr,
  output [31:0] io_coreRsp_bits_data,
  output [1:0]  io_coreRsp_bits_warpid,
  output [1:0]  io_coreRsp_bits_status,
  output        io_memRsp_ready,
  input         io_memRsp_valid,
  input  [31:0] io_memRsp_bits_d_addr,
  input  [31:0] io_memRsp_bits_d_data_0,
  input  [31:0] io_memRsp_bits_d_data_1,
  input  [31:0] io_memRsp_bits_d_data_2,
  input  [31:0] io_memRsp_bits_d_data_3,
  input  [31:0] io_memRsp_bits_d_data_4,
  input  [31:0] io_memRsp_bits_d_data_5,
  input  [31:0] io_memRsp_bits_d_data_6,
  input  [31:0] io_memRsp_bits_d_data_7,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [1:0]  io_memReq_bits_a_source,
  output [31:0] io_memReq_bits_a_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  tagAccess_clock; // @[ICache.scala 51:25]
  wire  tagAccess_reset; // @[ICache.scala 51:25]
  wire  tagAccess_io_r_req_valid; // @[ICache.scala 51:25]
  wire [4:0] tagAccess_io_r_req_bits_setIdx; // @[ICache.scala 51:25]
  wire [21:0] tagAccess_io_tagFromCore_st1; // @[ICache.scala 51:25]
  wire  tagAccess_io_coreReqReady; // @[ICache.scala 51:25]
  wire  tagAccess_io_w_req_valid; // @[ICache.scala 51:25]
  wire [4:0] tagAccess_io_w_req_bits_setIdx; // @[ICache.scala 51:25]
  wire [21:0] tagAccess_io_w_req_bits_data_0; // @[ICache.scala 51:25]
  wire [21:0] tagAccess_io_w_req_bits_data_1; // @[ICache.scala 51:25]
  wire [1:0] tagAccess_io_waymaskReplacement; // @[ICache.scala 51:25]
  wire [1:0] tagAccess_io_waymaskHit_st1; // @[ICache.scala 51:25]
  wire  tagAccess_io_hit_st1; // @[ICache.scala 51:25]
  wire  dataAccess_clock; // @[ICache.scala 52:26]
  wire  dataAccess_reset; // @[ICache.scala 52:26]
  wire  dataAccess_io_r_req_valid; // @[ICache.scala 52:26]
  wire [4:0] dataAccess_io_r_req_bits_setIdx; // @[ICache.scala 52:26]
  wire [255:0] dataAccess_io_r_resp_data_0; // @[ICache.scala 52:26]
  wire [255:0] dataAccess_io_r_resp_data_1; // @[ICache.scala 52:26]
  wire  dataAccess_io_w_req_valid; // @[ICache.scala 52:26]
  wire [4:0] dataAccess_io_w_req_bits_setIdx; // @[ICache.scala 52:26]
  wire [255:0] dataAccess_io_w_req_bits_data_0; // @[ICache.scala 52:26]
  wire [255:0] dataAccess_io_w_req_bits_data_1; // @[ICache.scala 52:26]
  wire [1:0] dataAccess_io_w_req_bits_waymask; // @[ICache.scala 52:26]
  wire  mshrAccess_clock; // @[ICache.scala 63:26]
  wire  mshrAccess_reset; // @[ICache.scala 63:26]
  wire  mshrAccess_io_missReq_ready; // @[ICache.scala 63:26]
  wire  mshrAccess_io_missReq_valid; // @[ICache.scala 63:26]
  wire [26:0] mshrAccess_io_missReq_bits_blockAddr; // @[ICache.scala 63:26]
  wire [1:0] mshrAccess_io_missReq_bits_targetInfo; // @[ICache.scala 63:26]
  wire  mshrAccess_io_missRspIn_ready; // @[ICache.scala 63:26]
  wire  mshrAccess_io_missRspIn_valid; // @[ICache.scala 63:26]
  wire [26:0] mshrAccess_io_missRspIn_bits_blockAddr; // @[ICache.scala 63:26]
  wire  mshrAccess_io_missRspOut_valid; // @[ICache.scala 63:26]
  wire [26:0] mshrAccess_io_missRspOut_bits_blockAddr; // @[ICache.scala 63:26]
  wire  mshrAccess_io_miss2mem_ready; // @[ICache.scala 63:26]
  wire  mshrAccess_io_miss2mem_valid; // @[ICache.scala 63:26]
  wire [26:0] mshrAccess_io_miss2mem_bits_blockAddr; // @[ICache.scala 63:26]
  wire [1:0] mshrAccess_io_miss2mem_bits_instrId; // @[ICache.scala 63:26]
  wire  memRsp_Q_clock; // @[ICache.scala 65:24]
  wire  memRsp_Q_reset; // @[ICache.scala 65:24]
  wire  memRsp_Q_io_enq_ready; // @[ICache.scala 65:24]
  wire  memRsp_Q_io_enq_valid; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_addr; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_0; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_1; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_2; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_3; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_4; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_5; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_6; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_7; // @[ICache.scala 65:24]
  wire  memRsp_Q_io_deq_ready; // @[ICache.scala 65:24]
  wire  memRsp_Q_io_deq_valid; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_addr; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_0; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_1; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_2; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_3; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_4; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_5; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_6; // @[ICache.scala 65:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_7; // @[ICache.scala 65:24]
  wire  _coreReqFire_st1_T = io_coreReq_ready & io_coreReq_valid; // @[Decoupled.scala 50:35]
  wire  ShouldFlushCoreRsp_st0 = io_coreReq_bits_warpid == io_externalFlushPipe_bits_warpid & io_externalFlushPipe_valid
    ; // @[ICache.scala 89:89]
  wire  _coreReqFire_st1_T_1 = ~ShouldFlushCoreRsp_st0; // @[ICache.scala 73:54]
  reg  coreReqFire_st1; // @[ICache.scala 73:32]
  reg [1:0] warpid_st1; // @[Reg.scala 16:16]
  wire  ShouldFlushCoreRsp_st1 = warpid_st1 == io_externalFlushPipe_bits_warpid & io_externalFlushPipe_valid; // @[ICache.scala 88:77]
  wire  _coreReqFire_st2_T = ~ShouldFlushCoreRsp_st1; // @[ICache.scala 74:52]
  reg  coreReqFire_st2; // @[ICache.scala 74:32]
  wire  cacheMiss_st1 = ~tagAccess_io_hit_st1 & coreReqFire_st1; // @[ICache.scala 76:45]
  wire  wayidx_hit_st1 = tagAccess_io_waymaskHit_st1[1]; // @[CircuitMath.scala 30:8]
  reg [1:0] warpid_st2; // @[ICache.scala 82:27]
  reg [31:0] addr_st1; // @[Reg.scala 16:16]
  reg [31:0] addr_st2; // @[ICache.scala 84:25]
  reg [31:0] pipeReqAddr_st1; // @[Reg.scala 16:16]
  wire [127:0] memRsp_QData_lo = {memRsp_Q_io_deq_bits_d_data_3,memRsp_Q_io_deq_bits_d_data_2,
    memRsp_Q_io_deq_bits_d_data_1,memRsp_Q_io_deq_bits_d_data_0}; // @[ICache.scala 104:53]
  wire [127:0] memRsp_QData_hi = {memRsp_Q_io_deq_bits_d_data_7,memRsp_Q_io_deq_bits_d_data_6,
    memRsp_Q_io_deq_bits_d_data_5,memRsp_Q_io_deq_bits_d_data_4}; // @[ICache.scala 104:53]
  wire [6:0] _mshrAccess_io_missReq_bits_targetInfo_T_1 = {warpid_st1,pipeReqAddr_st1[4:0]}; // @[Cat.scala 31:58]
  wire [511:0] _dataAccess_data_T = {dataAccess_io_r_resp_data_1,dataAccess_io_r_resp_data_0}; // @[ICache.scala 126:54]
  wire [255:0] dataAccess_data_0 = _dataAccess_data_T[255:0]; // @[ICache.scala 126:54]
  wire [255:0] dataAccess_data_1 = _dataAccess_data_T[511:256]; // @[ICache.scala 126:54]
  wire [2:0] blockOffset_sel_st1 = pipeReqAddr_st1[4:2]; // @[L1CacheParameters.scala 52:40]
  wire [7:0] _data_after_blockOffset_st1_T = {blockOffset_sel_st1, 5'h0}; // @[ICache.scala 130:85]
  wire [255:0] _GEN_4 = wayidx_hit_st1 ? dataAccess_data_1 : dataAccess_data_0; // @[ICache.scala 130:{61,61}]
  wire [255:0] _data_after_blockOffset_st1_T_1 = _GEN_4 >> _data_after_blockOffset_st1_T; // @[ICache.scala 130:61]
  reg [31:0] data_after_blockOffset_st2; // @[ICache.scala 132:43]
  reg  OrderViolation_st2; // @[ICache.scala 136:35]
  wire  _io_coreRsp_valid_T = ~OrderViolation_st2; // @[ICache.scala 137:42]
  reg  Status_st1_REG; // @[ICache.scala 152:31]
  wire  _Status_st1_T = mshrAccess_io_missReq_ready & mshrAccess_io_missReq_valid; // @[Decoupled.scala 50:35]
  wire  warpIdMatch2_st1 = warpid_st1 == warpid_st2; // @[ICache.scala 176:37]
  reg  cacheMiss_st2; // @[Reg.scala 16:16]
  reg [1:0] warpid_st3; // @[ICache.scala 172:27]
  wire  warpIdMatch3_st1 = warpid_st1 == warpid_st3; // @[ICache.scala 177:37]
  reg  cacheMiss_st3; // @[ICache.scala 174:30]
  reg  OrderViolation_st3; // @[ICache.scala 171:35]
  wire  OrderViolation_st1 = warpIdMatch2_st1 & cacheMiss_st2 & _io_coreRsp_valid_T | warpIdMatch3_st1 & cacheMiss_st3
     & ~OrderViolation_st3; // @[ICache.scala 179:84]
  wire  _Status_st1_T_3 = cacheMiss_st1 & ~_Status_st1_T | OrderViolation_st1; // @[ICache.scala 153:54]
  wire [1:0] _Status_st1_T_4 = {_Status_st1_T_3,cacheMiss_st1}; // @[Cat.scala 31:58]
  reg  Status_st2_REG; // @[ICache.scala 155:31]
  reg [1:0] Status_st2_REG_1; // @[ICache.scala 155:71]
  L1TagAccess tagAccess ( // @[ICache.scala 51:25]
    .clock(tagAccess_clock),
    .reset(tagAccess_reset),
    .io_r_req_valid(tagAccess_io_r_req_valid),
    .io_r_req_bits_setIdx(tagAccess_io_r_req_bits_setIdx),
    .io_tagFromCore_st1(tagAccess_io_tagFromCore_st1),
    .io_coreReqReady(tagAccess_io_coreReqReady),
    .io_w_req_valid(tagAccess_io_w_req_valid),
    .io_w_req_bits_setIdx(tagAccess_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(tagAccess_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(tagAccess_io_w_req_bits_data_1),
    .io_waymaskReplacement(tagAccess_io_waymaskReplacement),
    .io_waymaskHit_st1(tagAccess_io_waymaskHit_st1),
    .io_hit_st1(tagAccess_io_hit_st1)
  );
  SRAMTemplate_1 dataAccess ( // @[ICache.scala 52:26]
    .clock(dataAccess_clock),
    .reset(dataAccess_reset),
    .io_r_req_valid(dataAccess_io_r_req_valid),
    .io_r_req_bits_setIdx(dataAccess_io_r_req_bits_setIdx),
    .io_r_resp_data_0(dataAccess_io_r_resp_data_0),
    .io_r_resp_data_1(dataAccess_io_r_resp_data_1),
    .io_w_req_valid(dataAccess_io_w_req_valid),
    .io_w_req_bits_setIdx(dataAccess_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(dataAccess_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(dataAccess_io_w_req_bits_data_1),
    .io_w_req_bits_waymask(dataAccess_io_w_req_bits_waymask)
  );
  MSHR mshrAccess ( // @[ICache.scala 63:26]
    .clock(mshrAccess_clock),
    .reset(mshrAccess_reset),
    .io_missReq_ready(mshrAccess_io_missReq_ready),
    .io_missReq_valid(mshrAccess_io_missReq_valid),
    .io_missReq_bits_blockAddr(mshrAccess_io_missReq_bits_blockAddr),
    .io_missReq_bits_targetInfo(mshrAccess_io_missReq_bits_targetInfo),
    .io_missRspIn_ready(mshrAccess_io_missRspIn_ready),
    .io_missRspIn_valid(mshrAccess_io_missRspIn_valid),
    .io_missRspIn_bits_blockAddr(mshrAccess_io_missRspIn_bits_blockAddr),
    .io_missRspOut_valid(mshrAccess_io_missRspOut_valid),
    .io_missRspOut_bits_blockAddr(mshrAccess_io_missRspOut_bits_blockAddr),
    .io_miss2mem_ready(mshrAccess_io_miss2mem_ready),
    .io_miss2mem_valid(mshrAccess_io_miss2mem_valid),
    .io_miss2mem_bits_blockAddr(mshrAccess_io_miss2mem_bits_blockAddr),
    .io_miss2mem_bits_instrId(mshrAccess_io_miss2mem_bits_instrId)
  );
  Queue_49 memRsp_Q ( // @[ICache.scala 65:24]
    .clock(memRsp_Q_clock),
    .reset(memRsp_Q_reset),
    .io_enq_ready(memRsp_Q_io_enq_ready),
    .io_enq_valid(memRsp_Q_io_enq_valid),
    .io_enq_bits_d_addr(memRsp_Q_io_enq_bits_d_addr),
    .io_enq_bits_d_data_0(memRsp_Q_io_enq_bits_d_data_0),
    .io_enq_bits_d_data_1(memRsp_Q_io_enq_bits_d_data_1),
    .io_enq_bits_d_data_2(memRsp_Q_io_enq_bits_d_data_2),
    .io_enq_bits_d_data_3(memRsp_Q_io_enq_bits_d_data_3),
    .io_enq_bits_d_data_4(memRsp_Q_io_enq_bits_d_data_4),
    .io_enq_bits_d_data_5(memRsp_Q_io_enq_bits_d_data_5),
    .io_enq_bits_d_data_6(memRsp_Q_io_enq_bits_d_data_6),
    .io_enq_bits_d_data_7(memRsp_Q_io_enq_bits_d_data_7),
    .io_deq_ready(memRsp_Q_io_deq_ready),
    .io_deq_valid(memRsp_Q_io_deq_valid),
    .io_deq_bits_d_addr(memRsp_Q_io_deq_bits_d_addr),
    .io_deq_bits_d_data_0(memRsp_Q_io_deq_bits_d_data_0),
    .io_deq_bits_d_data_1(memRsp_Q_io_deq_bits_d_data_1),
    .io_deq_bits_d_data_2(memRsp_Q_io_deq_bits_d_data_2),
    .io_deq_bits_d_data_3(memRsp_Q_io_deq_bits_d_data_3),
    .io_deq_bits_d_data_4(memRsp_Q_io_deq_bits_d_data_4),
    .io_deq_bits_d_data_5(memRsp_Q_io_deq_bits_d_data_5),
    .io_deq_bits_d_data_6(memRsp_Q_io_deq_bits_d_data_6),
    .io_deq_bits_d_data_7(memRsp_Q_io_deq_bits_d_data_7)
  );
  assign io_coreReq_ready = 1'h1; // @[ICache.scala 165:20]
  assign io_coreRsp_valid = coreReqFire_st2 & ~OrderViolation_st2; // @[ICache.scala 137:39]
  assign io_coreRsp_bits_addr = addr_st2; // @[ICache.scala 145:24]
  assign io_coreRsp_bits_data = data_after_blockOffset_st2; // @[ICache.scala 138:24]
  assign io_coreRsp_bits_warpid = warpid_st2; // @[ICache.scala 139:26]
  assign io_coreRsp_bits_status = Status_st2_REG ? 2'h2 : Status_st2_REG_1; // @[ICache.scala 155:23]
  assign io_memRsp_ready = memRsp_Q_io_enq_ready; // @[ICache.scala 102:19]
  assign io_memReq_valid = mshrAccess_io_miss2mem_valid; // @[ICache.scala 158:19]
  assign io_memReq_bits_a_source = mshrAccess_io_miss2mem_bits_instrId; // @[ICache.scala 161:27]
  assign io_memReq_bits_a_addr = {mshrAccess_io_miss2mem_bits_blockAddr,5'h0}; // @[Cat.scala 31:58]
  assign tagAccess_clock = clock;
  assign tagAccess_reset = reset;
  assign tagAccess_io_r_req_valid = _coreReqFire_st1_T & _coreReqFire_st1_T_1; // @[ICache.scala 93:49]
  assign tagAccess_io_r_req_bits_setIdx = io_coreReq_bits_addr[9:5]; // @[L1CacheParameters.scala 45:9]
  assign tagAccess_io_tagFromCore_st1 = pipeReqAddr_st1[31:10]; // @[L1CacheParameters.scala 43:35]
  assign tagAccess_io_coreReqReady = io_coreReq_ready; // @[ICache.scala 96:29]
  assign tagAccess_io_w_req_valid = memRsp_Q_io_deq_ready & memRsp_Q_io_deq_valid; // @[Decoupled.scala 50:35]
  assign tagAccess_io_w_req_bits_setIdx = mshrAccess_io_missRspOut_bits_blockAddr[4:0]; // @[L1CacheParameters.scala 47:9]
  assign tagAccess_io_w_req_bits_data_0 = mshrAccess_io_missRspOut_bits_blockAddr[26:5]; // @[L1CacheParameters.scala 43:35]
  assign tagAccess_io_w_req_bits_data_1 = mshrAccess_io_missRspOut_bits_blockAddr[26:5]; // @[L1CacheParameters.scala 43:35]
  assign dataAccess_clock = clock;
  assign dataAccess_reset = reset;
  assign dataAccess_io_r_req_valid = _coreReqFire_st1_T & _coreReqFire_st1_T_1; // @[ICache.scala 124:50]
  assign dataAccess_io_r_req_bits_setIdx = io_coreReq_bits_addr[9:5]; // @[L1CacheParameters.scala 45:9]
  assign dataAccess_io_w_req_valid = memRsp_Q_io_deq_ready & memRsp_Q_io_deq_valid; // @[Decoupled.scala 50:35]
  assign dataAccess_io_w_req_bits_setIdx = mshrAccess_io_missRspOut_bits_blockAddr[4:0]; // @[L1CacheParameters.scala 47:9]
  assign dataAccess_io_w_req_bits_data_0 = {memRsp_QData_hi,memRsp_QData_lo}; // @[ICache.scala 104:53]
  assign dataAccess_io_w_req_bits_data_1 = {memRsp_QData_hi,memRsp_QData_lo}; // @[ICache.scala 104:53]
  assign dataAccess_io_w_req_bits_waymask = tagAccess_io_waymaskReplacement; // @[SRAMTemplate.scala 54:24]
  assign mshrAccess_clock = clock;
  assign mshrAccess_reset = reset;
  assign mshrAccess_io_missReq_valid = ~tagAccess_io_hit_st1 & coreReqFire_st1; // @[ICache.scala 76:45]
  assign mshrAccess_io_missReq_bits_blockAddr = pipeReqAddr_st1[31:5]; // @[L1CacheParameters.scala 55:41]
  assign mshrAccess_io_missReq_bits_targetInfo = _mshrAccess_io_missReq_bits_targetInfo_T_1[1:0]; // @[ICache.scala 109:41]
  assign mshrAccess_io_missRspIn_valid = memRsp_Q_io_deq_valid; // @[ICache.scala 113:33]
  assign mshrAccess_io_missRspIn_bits_blockAddr = memRsp_Q_io_deq_bits_d_addr[31:5]; // @[L1CacheParameters.scala 55:41]
  assign mshrAccess_io_miss2mem_ready = io_memReq_ready; // @[ICache.scala 159:32]
  assign memRsp_Q_clock = clock;
  assign memRsp_Q_reset = reset;
  assign memRsp_Q_io_enq_valid = io_memRsp_valid; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_addr = io_memRsp_bits_d_addr; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_0 = io_memRsp_bits_d_data_0; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_1 = io_memRsp_bits_d_data_1; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_2 = io_memRsp_bits_d_data_2; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_3 = io_memRsp_bits_d_data_3; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_4 = io_memRsp_bits_d_data_4; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_5 = io_memRsp_bits_d_data_5; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_6 = io_memRsp_bits_d_data_6; // @[ICache.scala 102:19]
  assign memRsp_Q_io_enq_bits_d_data_7 = io_memRsp_bits_d_data_7; // @[ICache.scala 102:19]
  assign memRsp_Q_io_deq_ready = mshrAccess_io_missRspIn_ready; // @[ICache.scala 112:25]
  always @(posedge clock) begin
    coreReqFire_st1 <= _coreReqFire_st1_T & ~ShouldFlushCoreRsp_st0; // @[ICache.scala 73:51]
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      warpid_st1 <= io_coreReq_bits_warpid; // @[Reg.scala 17:22]
    end
    coreReqFire_st2 <= coreReqFire_st1 & ~ShouldFlushCoreRsp_st1; // @[ICache.scala 74:49]
    warpid_st2 <= warpid_st1; // @[ICache.scala 82:27]
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      addr_st1 <= io_coreReq_bits_addr; // @[Reg.scala 17:22]
    end
    addr_st2 <= addr_st1; // @[ICache.scala 84:25]
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      pipeReqAddr_st1 <= io_coreReq_bits_addr; // @[Reg.scala 17:22]
    end
    data_after_blockOffset_st2 <= _data_after_blockOffset_st1_T_1[31:0]; // @[ICache.scala 130:91]
    OrderViolation_st2 <= warpIdMatch2_st1 & cacheMiss_st2 & _io_coreRsp_valid_T | warpIdMatch3_st1 & cacheMiss_st3 & ~
      OrderViolation_st3; // @[ICache.scala 179:84]
    Status_st1_REG <= io_coreReq_bits_warpid == io_externalFlushPipe_bits_warpid & io_externalFlushPipe_valid; // @[ICache.scala 89:89]
    if (_coreReqFire_st2_T) begin // @[Reg.scala 17:18]
      cacheMiss_st2 <= cacheMiss_st1; // @[Reg.scala 17:22]
    end
    warpid_st3 <= warpid_st2; // @[ICache.scala 172:27]
    cacheMiss_st3 <= cacheMiss_st2; // @[ICache.scala 174:30]
    OrderViolation_st3 <= OrderViolation_st2; // @[ICache.scala 171:35]
    Status_st2_REG <= warpid_st1 == io_externalFlushPipe_bits_warpid & io_externalFlushPipe_valid; // @[ICache.scala 88:77]
    if (Status_st1_REG) begin // @[ICache.scala 152:23]
      Status_st2_REG_1 <= 2'h2;
    end else begin
      Status_st2_REG_1 <= _Status_st1_T_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  coreReqFire_st1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  warpid_st1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  coreReqFire_st2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  warpid_st2 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  addr_st1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  addr_st2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  pipeReqAddr_st1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  data_after_blockOffset_st2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  OrderViolation_st2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  Status_st1_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  cacheMiss_st2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  warpid_st3 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  cacheMiss_st3 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  OrderViolation_st3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  Status_st2_REG = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  Status_st2_REG_1 = _RAND_15[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BankConflictArbiter(
  input        clock,
  input        reset,
  input        io_coreReqArb_isWrite,
  input        io_coreReqArb_enable,
  input        io_coreReqArb_perLaneAddr_0_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_0_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_0_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_1_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_1_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_1_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_2_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_2_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_2_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_3_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_3_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_3_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_4_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_4_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_4_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_5_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_5_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_5_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_6_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_6_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_6_wordOffset1H,
  input        io_coreReqArb_perLaneAddr_7_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_7_blockOffset,
  input  [3:0] io_coreReqArb_perLaneAddr_7_wordOffset1H,
  output [7:0] io_dataCrsbarSel1H_0,
  output [7:0] io_dataCrsbarSel1H_1,
  output [7:0] io_dataCrsbarSel1H_2,
  output [7:0] io_dataCrsbarSel1H_3,
  output [7:0] io_dataCrsbarSel1H_4,
  output [7:0] io_dataCrsbarSel1H_5,
  output [7:0] io_dataCrsbarSel1H_6,
  output [7:0] io_dataCrsbarSel1H_7,
  output [3:0] io_addrCrsbarOut_0_wordOffset1H,
  output [3:0] io_addrCrsbarOut_1_wordOffset1H,
  output [3:0] io_addrCrsbarOut_2_wordOffset1H,
  output [3:0] io_addrCrsbarOut_3_wordOffset1H,
  output [3:0] io_addrCrsbarOut_4_wordOffset1H,
  output [3:0] io_addrCrsbarOut_5_wordOffset1H,
  output [3:0] io_addrCrsbarOut_6_wordOffset1H,
  output [3:0] io_addrCrsbarOut_7_wordOffset1H,
  output       io_dataArrayEn_0,
  output       io_dataArrayEn_1,
  output       io_dataArrayEn_2,
  output       io_dataArrayEn_3,
  output       io_dataArrayEn_4,
  output       io_dataArrayEn_5,
  output       io_dataArrayEn_6,
  output       io_dataArrayEn_7,
  output       io_activeLane_0,
  output       io_activeLane_1,
  output       io_activeLane_2,
  output       io_activeLane_3,
  output       io_activeLane_4,
  output       io_activeLane_5,
  output       io_activeLane_6,
  output       io_activeLane_7,
  output       io_bankConflict
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  reg  bankConflict_reg; // @[BankConflictArbiter.scala 105:33]
  reg  conflictReqIsW_reg; // @[BankConflictArbiter.scala 106:31]
  reg  perLaneConflictReq_reg_0_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_0_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_0_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_1_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_1_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_1_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_2_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_2_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_2_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_3_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_3_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_3_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_4_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_4_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_4_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_5_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_5_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_5_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_6_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_6_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_6_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  reg  perLaneConflictReq_reg_7_activeMask; // @[BankConflictArbiter.scala 108:35]
  reg [2:0] perLaneConflictReq_reg_7_bankIdx; // @[BankConflictArbiter.scala 108:35]
  reg [3:0] perLaneConflictReq_reg_7_AddrBundle_wordOffset1H; // @[BankConflictArbiter.scala 108:35]
  wire  isWrite = bankConflict_reg ? conflictReqIsW_reg : io_coreReqArb_isWrite; // @[BankConflictArbiter.scala 123:26]
  wire [2:0] perLaneConflictReq_0_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_0_bankIdx :
    io_coreReqArb_perLaneAddr_0_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_0 = 8'h1 << perLaneConflictReq_0_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_0_activeMask = bankConflict_reg ? perLaneConflictReq_reg_0_activeMask :
    io_coreReqArb_perLaneAddr_0_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_0_T_1 = perLaneConflictReq_0_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_0 = bankIdx1H_0 & _bankIdxMasked_0_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_1_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_1_bankIdx :
    io_coreReqArb_perLaneAddr_1_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_1 = 8'h1 << perLaneConflictReq_1_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_1_activeMask = bankConflict_reg ? perLaneConflictReq_reg_1_activeMask :
    io_coreReqArb_perLaneAddr_1_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_1_T_1 = perLaneConflictReq_1_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_1 = bankIdx1H_1 & _bankIdxMasked_1_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_2_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_2_bankIdx :
    io_coreReqArb_perLaneAddr_2_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_2 = 8'h1 << perLaneConflictReq_2_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_2_activeMask = bankConflict_reg ? perLaneConflictReq_reg_2_activeMask :
    io_coreReqArb_perLaneAddr_2_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_2_T_1 = perLaneConflictReq_2_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_2 = bankIdx1H_2 & _bankIdxMasked_2_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_3_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_3_bankIdx :
    io_coreReqArb_perLaneAddr_3_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_3 = 8'h1 << perLaneConflictReq_3_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_3_activeMask = bankConflict_reg ? perLaneConflictReq_reg_3_activeMask :
    io_coreReqArb_perLaneAddr_3_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_3_T_1 = perLaneConflictReq_3_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_3 = bankIdx1H_3 & _bankIdxMasked_3_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_4_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_4_bankIdx :
    io_coreReqArb_perLaneAddr_4_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_4 = 8'h1 << perLaneConflictReq_4_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_4_activeMask = bankConflict_reg ? perLaneConflictReq_reg_4_activeMask :
    io_coreReqArb_perLaneAddr_4_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_4_T_1 = perLaneConflictReq_4_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_4 = bankIdx1H_4 & _bankIdxMasked_4_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_5_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_5_bankIdx :
    io_coreReqArb_perLaneAddr_5_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_5 = 8'h1 << perLaneConflictReq_5_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_5_activeMask = bankConflict_reg ? perLaneConflictReq_reg_5_activeMask :
    io_coreReqArb_perLaneAddr_5_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_5_T_1 = perLaneConflictReq_5_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_5 = bankIdx1H_5 & _bankIdxMasked_5_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_6_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_6_bankIdx :
    io_coreReqArb_perLaneAddr_6_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_6 = 8'h1 << perLaneConflictReq_6_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_6_activeMask = bankConflict_reg ? perLaneConflictReq_reg_6_activeMask :
    io_coreReqArb_perLaneAddr_6_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_6_T_1 = perLaneConflictReq_6_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_6 = bankIdx1H_6 & _bankIdxMasked_6_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [2:0] perLaneConflictReq_7_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_7_bankIdx :
    io_coreReqArb_perLaneAddr_7_blockOffset; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] bankIdx1H_7 = 8'h1 << perLaneConflictReq_7_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_7_activeMask = bankConflict_reg ? perLaneConflictReq_reg_7_activeMask :
    io_coreReqArb_perLaneAddr_7_activeMask; // @[BankConflictArbiter.scala 159:28]
  wire [7:0] _bankIdxMasked_7_T_1 = perLaneConflictReq_7_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_7 = bankIdx1H_7 & _bankIdxMasked_7_T_1; // @[BankConflictArbiter.scala 131:38]
  wire [7:0] _perBankReq_Bin_0_T_8 = {bankIdxMasked_0[0],bankIdxMasked_1[0],bankIdxMasked_2[0],bankIdxMasked_3[0],
    bankIdxMasked_4[0],bankIdxMasked_5[0],bankIdxMasked_6[0],bankIdxMasked_7[0]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_17 = {{4'd0}, _perBankReq_Bin_0_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_12 = _GEN_17 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_14 = {_perBankReq_Bin_0_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_0_T_16 = _perBankReq_Bin_0_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_0_T_17 = _perBankReq_Bin_0_T_12 | _perBankReq_Bin_0_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_18 = {{2'd0}, _perBankReq_Bin_0_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_22 = _GEN_18 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_24 = {_perBankReq_Bin_0_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_0_T_26 = _perBankReq_Bin_0_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_0_T_27 = _perBankReq_Bin_0_T_22 | _perBankReq_Bin_0_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_19 = {{1'd0}, _perBankReq_Bin_0_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_32 = _GEN_19 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_34 = {_perBankReq_Bin_0_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_0_T_36 = _perBankReq_Bin_0_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_0 = _perBankReq_Bin_0_T_32 | _perBankReq_Bin_0_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_0_T_8 = perBankReq_Bin_0[0] + perBankReq_Bin_0[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_0_T_10 = perBankReq_Bin_0[2] + perBankReq_Bin_0[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_0_T_12 = _perBankReqCount_0_T_8 + _perBankReqCount_0_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_0_T_14 = perBankReq_Bin_0[4] + perBankReq_Bin_0[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_0_T_16 = perBankReq_Bin_0[6] + perBankReq_Bin_0[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_0_T_18 = _perBankReqCount_0_T_14 + _perBankReqCount_0_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_0_T_20 = _perBankReqCount_0_T_12 + _perBankReqCount_0_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_1_T_8 = {bankIdxMasked_0[1],bankIdxMasked_1[1],bankIdxMasked_2[1],bankIdxMasked_3[1],
    bankIdxMasked_4[1],bankIdxMasked_5[1],bankIdxMasked_6[1],bankIdxMasked_7[1]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_20 = {{4'd0}, _perBankReq_Bin_1_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_12 = _GEN_20 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_14 = {_perBankReq_Bin_1_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_1_T_16 = _perBankReq_Bin_1_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_1_T_17 = _perBankReq_Bin_1_T_12 | _perBankReq_Bin_1_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_21 = {{2'd0}, _perBankReq_Bin_1_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_22 = _GEN_21 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_24 = {_perBankReq_Bin_1_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_1_T_26 = _perBankReq_Bin_1_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_1_T_27 = _perBankReq_Bin_1_T_22 | _perBankReq_Bin_1_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_22 = {{1'd0}, _perBankReq_Bin_1_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_32 = _GEN_22 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_34 = {_perBankReq_Bin_1_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_1_T_36 = _perBankReq_Bin_1_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_1 = _perBankReq_Bin_1_T_32 | _perBankReq_Bin_1_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_1_T_8 = perBankReq_Bin_1[0] + perBankReq_Bin_1[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_1_T_10 = perBankReq_Bin_1[2] + perBankReq_Bin_1[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_1_T_12 = _perBankReqCount_1_T_8 + _perBankReqCount_1_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_1_T_14 = perBankReq_Bin_1[4] + perBankReq_Bin_1[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_1_T_16 = perBankReq_Bin_1[6] + perBankReq_Bin_1[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_1_T_18 = _perBankReqCount_1_T_14 + _perBankReqCount_1_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_1_T_20 = _perBankReqCount_1_T_12 + _perBankReqCount_1_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_2_T_8 = {bankIdxMasked_0[2],bankIdxMasked_1[2],bankIdxMasked_2[2],bankIdxMasked_3[2],
    bankIdxMasked_4[2],bankIdxMasked_5[2],bankIdxMasked_6[2],bankIdxMasked_7[2]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_23 = {{4'd0}, _perBankReq_Bin_2_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_12 = _GEN_23 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_14 = {_perBankReq_Bin_2_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_2_T_16 = _perBankReq_Bin_2_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_2_T_17 = _perBankReq_Bin_2_T_12 | _perBankReq_Bin_2_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_24 = {{2'd0}, _perBankReq_Bin_2_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_22 = _GEN_24 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_24 = {_perBankReq_Bin_2_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_2_T_26 = _perBankReq_Bin_2_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_2_T_27 = _perBankReq_Bin_2_T_22 | _perBankReq_Bin_2_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_25 = {{1'd0}, _perBankReq_Bin_2_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_32 = _GEN_25 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_34 = {_perBankReq_Bin_2_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_2_T_36 = _perBankReq_Bin_2_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_2 = _perBankReq_Bin_2_T_32 | _perBankReq_Bin_2_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_2_T_8 = perBankReq_Bin_2[0] + perBankReq_Bin_2[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_2_T_10 = perBankReq_Bin_2[2] + perBankReq_Bin_2[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_2_T_12 = _perBankReqCount_2_T_8 + _perBankReqCount_2_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_2_T_14 = perBankReq_Bin_2[4] + perBankReq_Bin_2[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_2_T_16 = perBankReq_Bin_2[6] + perBankReq_Bin_2[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_2_T_18 = _perBankReqCount_2_T_14 + _perBankReqCount_2_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_2_T_20 = _perBankReqCount_2_T_12 + _perBankReqCount_2_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_3_T_8 = {bankIdxMasked_0[3],bankIdxMasked_1[3],bankIdxMasked_2[3],bankIdxMasked_3[3],
    bankIdxMasked_4[3],bankIdxMasked_5[3],bankIdxMasked_6[3],bankIdxMasked_7[3]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_26 = {{4'd0}, _perBankReq_Bin_3_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_12 = _GEN_26 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_14 = {_perBankReq_Bin_3_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_3_T_16 = _perBankReq_Bin_3_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_3_T_17 = _perBankReq_Bin_3_T_12 | _perBankReq_Bin_3_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_27 = {{2'd0}, _perBankReq_Bin_3_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_22 = _GEN_27 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_24 = {_perBankReq_Bin_3_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_3_T_26 = _perBankReq_Bin_3_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_3_T_27 = _perBankReq_Bin_3_T_22 | _perBankReq_Bin_3_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_28 = {{1'd0}, _perBankReq_Bin_3_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_32 = _GEN_28 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_34 = {_perBankReq_Bin_3_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_3_T_36 = _perBankReq_Bin_3_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_3 = _perBankReq_Bin_3_T_32 | _perBankReq_Bin_3_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_3_T_8 = perBankReq_Bin_3[0] + perBankReq_Bin_3[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_3_T_10 = perBankReq_Bin_3[2] + perBankReq_Bin_3[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_3_T_12 = _perBankReqCount_3_T_8 + _perBankReqCount_3_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_3_T_14 = perBankReq_Bin_3[4] + perBankReq_Bin_3[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_3_T_16 = perBankReq_Bin_3[6] + perBankReq_Bin_3[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_3_T_18 = _perBankReqCount_3_T_14 + _perBankReqCount_3_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_3_T_20 = _perBankReqCount_3_T_12 + _perBankReqCount_3_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_4_T_8 = {bankIdxMasked_0[4],bankIdxMasked_1[4],bankIdxMasked_2[4],bankIdxMasked_3[4],
    bankIdxMasked_4[4],bankIdxMasked_5[4],bankIdxMasked_6[4],bankIdxMasked_7[4]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_29 = {{4'd0}, _perBankReq_Bin_4_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_12 = _GEN_29 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_14 = {_perBankReq_Bin_4_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_4_T_16 = _perBankReq_Bin_4_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_4_T_17 = _perBankReq_Bin_4_T_12 | _perBankReq_Bin_4_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_30 = {{2'd0}, _perBankReq_Bin_4_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_22 = _GEN_30 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_24 = {_perBankReq_Bin_4_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_4_T_26 = _perBankReq_Bin_4_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_4_T_27 = _perBankReq_Bin_4_T_22 | _perBankReq_Bin_4_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_31 = {{1'd0}, _perBankReq_Bin_4_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_32 = _GEN_31 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_34 = {_perBankReq_Bin_4_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_4_T_36 = _perBankReq_Bin_4_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_4 = _perBankReq_Bin_4_T_32 | _perBankReq_Bin_4_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_4_T_8 = perBankReq_Bin_4[0] + perBankReq_Bin_4[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_4_T_10 = perBankReq_Bin_4[2] + perBankReq_Bin_4[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_4_T_12 = _perBankReqCount_4_T_8 + _perBankReqCount_4_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_4_T_14 = perBankReq_Bin_4[4] + perBankReq_Bin_4[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_4_T_16 = perBankReq_Bin_4[6] + perBankReq_Bin_4[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_4_T_18 = _perBankReqCount_4_T_14 + _perBankReqCount_4_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_4_T_20 = _perBankReqCount_4_T_12 + _perBankReqCount_4_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_5_T_8 = {bankIdxMasked_0[5],bankIdxMasked_1[5],bankIdxMasked_2[5],bankIdxMasked_3[5],
    bankIdxMasked_4[5],bankIdxMasked_5[5],bankIdxMasked_6[5],bankIdxMasked_7[5]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_32 = {{4'd0}, _perBankReq_Bin_5_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_12 = _GEN_32 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_14 = {_perBankReq_Bin_5_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_5_T_16 = _perBankReq_Bin_5_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_5_T_17 = _perBankReq_Bin_5_T_12 | _perBankReq_Bin_5_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_33 = {{2'd0}, _perBankReq_Bin_5_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_22 = _GEN_33 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_24 = {_perBankReq_Bin_5_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_5_T_26 = _perBankReq_Bin_5_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_5_T_27 = _perBankReq_Bin_5_T_22 | _perBankReq_Bin_5_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_34 = {{1'd0}, _perBankReq_Bin_5_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_32 = _GEN_34 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_34 = {_perBankReq_Bin_5_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_5_T_36 = _perBankReq_Bin_5_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_5 = _perBankReq_Bin_5_T_32 | _perBankReq_Bin_5_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_5_T_8 = perBankReq_Bin_5[0] + perBankReq_Bin_5[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_5_T_10 = perBankReq_Bin_5[2] + perBankReq_Bin_5[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_5_T_12 = _perBankReqCount_5_T_8 + _perBankReqCount_5_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_5_T_14 = perBankReq_Bin_5[4] + perBankReq_Bin_5[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_5_T_16 = perBankReq_Bin_5[6] + perBankReq_Bin_5[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_5_T_18 = _perBankReqCount_5_T_14 + _perBankReqCount_5_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_5_T_20 = _perBankReqCount_5_T_12 + _perBankReqCount_5_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_6_T_8 = {bankIdxMasked_0[6],bankIdxMasked_1[6],bankIdxMasked_2[6],bankIdxMasked_3[6],
    bankIdxMasked_4[6],bankIdxMasked_5[6],bankIdxMasked_6[6],bankIdxMasked_7[6]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_35 = {{4'd0}, _perBankReq_Bin_6_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_12 = _GEN_35 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_14 = {_perBankReq_Bin_6_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_6_T_16 = _perBankReq_Bin_6_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_6_T_17 = _perBankReq_Bin_6_T_12 | _perBankReq_Bin_6_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_36 = {{2'd0}, _perBankReq_Bin_6_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_22 = _GEN_36 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_24 = {_perBankReq_Bin_6_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_6_T_26 = _perBankReq_Bin_6_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_6_T_27 = _perBankReq_Bin_6_T_22 | _perBankReq_Bin_6_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_37 = {{1'd0}, _perBankReq_Bin_6_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_32 = _GEN_37 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_34 = {_perBankReq_Bin_6_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_6_T_36 = _perBankReq_Bin_6_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_6 = _perBankReq_Bin_6_T_32 | _perBankReq_Bin_6_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_6_T_8 = perBankReq_Bin_6[0] + perBankReq_Bin_6[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_6_T_10 = perBankReq_Bin_6[2] + perBankReq_Bin_6[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_6_T_12 = _perBankReqCount_6_T_8 + _perBankReqCount_6_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_6_T_14 = perBankReq_Bin_6[4] + perBankReq_Bin_6[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_6_T_16 = perBankReq_Bin_6[6] + perBankReq_Bin_6[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_6_T_18 = _perBankReqCount_6_T_14 + _perBankReqCount_6_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_6_T_20 = _perBankReqCount_6_T_12 + _perBankReqCount_6_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_7_T_8 = {bankIdxMasked_0[7],bankIdxMasked_1[7],bankIdxMasked_2[7],bankIdxMasked_3[7],
    bankIdxMasked_4[7],bankIdxMasked_5[7],bankIdxMasked_6[7],bankIdxMasked_7[7]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_38 = {{4'd0}, _perBankReq_Bin_7_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_12 = _GEN_38 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_14 = {_perBankReq_Bin_7_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_7_T_16 = _perBankReq_Bin_7_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_7_T_17 = _perBankReq_Bin_7_T_12 | _perBankReq_Bin_7_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_39 = {{2'd0}, _perBankReq_Bin_7_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_22 = _GEN_39 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_24 = {_perBankReq_Bin_7_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_7_T_26 = _perBankReq_Bin_7_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_7_T_27 = _perBankReq_Bin_7_T_22 | _perBankReq_Bin_7_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_40 = {{1'd0}, _perBankReq_Bin_7_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_32 = _GEN_40 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_34 = {_perBankReq_Bin_7_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_7_T_36 = _perBankReq_Bin_7_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_7 = _perBankReq_Bin_7_T_32 | _perBankReq_Bin_7_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_7_T_8 = perBankReq_Bin_7[0] + perBankReq_Bin_7[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_7_T_10 = perBankReq_Bin_7[2] + perBankReq_Bin_7[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_7_T_12 = _perBankReqCount_7_T_8 + _perBankReqCount_7_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_7_T_14 = perBankReq_Bin_7[4] + perBankReq_Bin_7[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_7_T_16 = perBankReq_Bin_7[6] + perBankReq_Bin_7[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_7_T_18 = _perBankReqCount_7_T_14 + _perBankReqCount_7_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_7_T_20 = _perBankReqCount_7_T_12 + _perBankReqCount_7_T_18; // @[Bitwise.scala 48:55]
  wire [2:0] perBankReqCount_0 = _perBankReqCount_0_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_0 = perBankReqCount_0 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_1 = _perBankReqCount_1_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_1 = perBankReqCount_1 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_2 = _perBankReqCount_2_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_2 = perBankReqCount_2 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_3 = _perBankReqCount_3_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_3 = perBankReqCount_3 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_4 = _perBankReqCount_4_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_4 = perBankReqCount_4 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_5 = _perBankReqCount_5_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_5 = perBankReqCount_5 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_6 = _perBankReqCount_6_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_6 = perBankReqCount_6 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [2:0] perBankReqCount_7 = _perBankReqCount_7_T_20[2:0]; // @[BankConflictArbiter.scala 133:29 136:24]
  wire  perBankReqConflict_7 = perBankReqCount_7 > 3'h1; // @[BankConflictArbiter.scala 147:46]
  wire [7:0] _bankConflict_T = {perBankReqConflict_0,perBankReqConflict_1,perBankReqConflict_2,perBankReqConflict_3,
    perBankReqConflict_4,perBankReqConflict_5,perBankReqConflict_6,perBankReqConflict_7}; // @[Cat.scala 31:58]
  wire  bankConflict = |_bankConflict_T & (io_coreReqArb_enable | bankConflict_reg); // @[BankConflictArbiter.scala 148:47]
  wire [7:0] _T_16 = perBankReq_Bin_0[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_17 = perBankReq_Bin_0[6] ? 8'h40 : _T_16; // @[Mux.scala 47:70]
  wire [7:0] _T_18 = perBankReq_Bin_0[5] ? 8'h20 : _T_17; // @[Mux.scala 47:70]
  wire [7:0] _T_19 = perBankReq_Bin_0[4] ? 8'h10 : _T_18; // @[Mux.scala 47:70]
  wire [7:0] _T_20 = perBankReq_Bin_0[3] ? 8'h8 : _T_19; // @[Mux.scala 47:70]
  wire [7:0] _T_21 = perBankReq_Bin_0[2] ? 8'h4 : _T_20; // @[Mux.scala 47:70]
  wire [7:0] _T_22 = perBankReq_Bin_0[1] ? 8'h2 : _T_21; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_0 = perBankReq_Bin_0[0] ? 8'h1 : _T_22; // @[Mux.scala 47:70]
  wire [7:0] _T_32 = perBankReq_Bin_1[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_33 = perBankReq_Bin_1[6] ? 8'h40 : _T_32; // @[Mux.scala 47:70]
  wire [7:0] _T_34 = perBankReq_Bin_1[5] ? 8'h20 : _T_33; // @[Mux.scala 47:70]
  wire [7:0] _T_35 = perBankReq_Bin_1[4] ? 8'h10 : _T_34; // @[Mux.scala 47:70]
  wire [7:0] _T_36 = perBankReq_Bin_1[3] ? 8'h8 : _T_35; // @[Mux.scala 47:70]
  wire [7:0] _T_37 = perBankReq_Bin_1[2] ? 8'h4 : _T_36; // @[Mux.scala 47:70]
  wire [7:0] _T_38 = perBankReq_Bin_1[1] ? 8'h2 : _T_37; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_1 = perBankReq_Bin_1[0] ? 8'h1 : _T_38; // @[Mux.scala 47:70]
  wire [7:0] _T_48 = perBankReq_Bin_2[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_49 = perBankReq_Bin_2[6] ? 8'h40 : _T_48; // @[Mux.scala 47:70]
  wire [7:0] _T_50 = perBankReq_Bin_2[5] ? 8'h20 : _T_49; // @[Mux.scala 47:70]
  wire [7:0] _T_51 = perBankReq_Bin_2[4] ? 8'h10 : _T_50; // @[Mux.scala 47:70]
  wire [7:0] _T_52 = perBankReq_Bin_2[3] ? 8'h8 : _T_51; // @[Mux.scala 47:70]
  wire [7:0] _T_53 = perBankReq_Bin_2[2] ? 8'h4 : _T_52; // @[Mux.scala 47:70]
  wire [7:0] _T_54 = perBankReq_Bin_2[1] ? 8'h2 : _T_53; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_2 = perBankReq_Bin_2[0] ? 8'h1 : _T_54; // @[Mux.scala 47:70]
  wire [7:0] _T_64 = perBankReq_Bin_3[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_65 = perBankReq_Bin_3[6] ? 8'h40 : _T_64; // @[Mux.scala 47:70]
  wire [7:0] _T_66 = perBankReq_Bin_3[5] ? 8'h20 : _T_65; // @[Mux.scala 47:70]
  wire [7:0] _T_67 = perBankReq_Bin_3[4] ? 8'h10 : _T_66; // @[Mux.scala 47:70]
  wire [7:0] _T_68 = perBankReq_Bin_3[3] ? 8'h8 : _T_67; // @[Mux.scala 47:70]
  wire [7:0] _T_69 = perBankReq_Bin_3[2] ? 8'h4 : _T_68; // @[Mux.scala 47:70]
  wire [7:0] _T_70 = perBankReq_Bin_3[1] ? 8'h2 : _T_69; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_3 = perBankReq_Bin_3[0] ? 8'h1 : _T_70; // @[Mux.scala 47:70]
  wire [7:0] _T_80 = perBankReq_Bin_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_81 = perBankReq_Bin_4[6] ? 8'h40 : _T_80; // @[Mux.scala 47:70]
  wire [7:0] _T_82 = perBankReq_Bin_4[5] ? 8'h20 : _T_81; // @[Mux.scala 47:70]
  wire [7:0] _T_83 = perBankReq_Bin_4[4] ? 8'h10 : _T_82; // @[Mux.scala 47:70]
  wire [7:0] _T_84 = perBankReq_Bin_4[3] ? 8'h8 : _T_83; // @[Mux.scala 47:70]
  wire [7:0] _T_85 = perBankReq_Bin_4[2] ? 8'h4 : _T_84; // @[Mux.scala 47:70]
  wire [7:0] _T_86 = perBankReq_Bin_4[1] ? 8'h2 : _T_85; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_4 = perBankReq_Bin_4[0] ? 8'h1 : _T_86; // @[Mux.scala 47:70]
  wire [7:0] _T_96 = perBankReq_Bin_5[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_97 = perBankReq_Bin_5[6] ? 8'h40 : _T_96; // @[Mux.scala 47:70]
  wire [7:0] _T_98 = perBankReq_Bin_5[5] ? 8'h20 : _T_97; // @[Mux.scala 47:70]
  wire [7:0] _T_99 = perBankReq_Bin_5[4] ? 8'h10 : _T_98; // @[Mux.scala 47:70]
  wire [7:0] _T_100 = perBankReq_Bin_5[3] ? 8'h8 : _T_99; // @[Mux.scala 47:70]
  wire [7:0] _T_101 = perBankReq_Bin_5[2] ? 8'h4 : _T_100; // @[Mux.scala 47:70]
  wire [7:0] _T_102 = perBankReq_Bin_5[1] ? 8'h2 : _T_101; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_5 = perBankReq_Bin_5[0] ? 8'h1 : _T_102; // @[Mux.scala 47:70]
  wire [7:0] _T_112 = perBankReq_Bin_6[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_113 = perBankReq_Bin_6[6] ? 8'h40 : _T_112; // @[Mux.scala 47:70]
  wire [7:0] _T_114 = perBankReq_Bin_6[5] ? 8'h20 : _T_113; // @[Mux.scala 47:70]
  wire [7:0] _T_115 = perBankReq_Bin_6[4] ? 8'h10 : _T_114; // @[Mux.scala 47:70]
  wire [7:0] _T_116 = perBankReq_Bin_6[3] ? 8'h8 : _T_115; // @[Mux.scala 47:70]
  wire [7:0] _T_117 = perBankReq_Bin_6[2] ? 8'h4 : _T_116; // @[Mux.scala 47:70]
  wire [7:0] _T_118 = perBankReq_Bin_6[1] ? 8'h2 : _T_117; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_6 = perBankReq_Bin_6[0] ? 8'h1 : _T_118; // @[Mux.scala 47:70]
  wire [7:0] _T_128 = perBankReq_Bin_7[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_129 = perBankReq_Bin_7[6] ? 8'h40 : _T_128; // @[Mux.scala 47:70]
  wire [7:0] _T_130 = perBankReq_Bin_7[5] ? 8'h20 : _T_129; // @[Mux.scala 47:70]
  wire [7:0] _T_131 = perBankReq_Bin_7[4] ? 8'h10 : _T_130; // @[Mux.scala 47:70]
  wire [7:0] _T_132 = perBankReq_Bin_7[3] ? 8'h8 : _T_131; // @[Mux.scala 47:70]
  wire [7:0] _T_133 = perBankReq_Bin_7[2] ? 8'h4 : _T_132; // @[Mux.scala 47:70]
  wire [7:0] _T_134 = perBankReq_Bin_7[1] ? 8'h2 : _T_133; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_7 = perBankReq_Bin_7[0] ? 8'h1 : _T_134; // @[Mux.scala 47:70]
  wire [7:0] _ActiveLaneWhenConflict1H_0_T_8 = {perBankActiveLaneWhenConflict1H_0[0],perBankActiveLaneWhenConflict1H_1[0
    ],perBankActiveLaneWhenConflict1H_2[0],perBankActiveLaneWhenConflict1H_3[0],perBankActiveLaneWhenConflict1H_4[0],
    perBankActiveLaneWhenConflict1H_5[0],perBankActiveLaneWhenConflict1H_6[0],perBankActiveLaneWhenConflict1H_7[0]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_0 = |_ActiveLaneWhenConflict1H_0_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_1_T_8 = {perBankActiveLaneWhenConflict1H_0[1],perBankActiveLaneWhenConflict1H_1[1
    ],perBankActiveLaneWhenConflict1H_2[1],perBankActiveLaneWhenConflict1H_3[1],perBankActiveLaneWhenConflict1H_4[1],
    perBankActiveLaneWhenConflict1H_5[1],perBankActiveLaneWhenConflict1H_6[1],perBankActiveLaneWhenConflict1H_7[1]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_1 = |_ActiveLaneWhenConflict1H_1_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_2_T_8 = {perBankActiveLaneWhenConflict1H_0[2],perBankActiveLaneWhenConflict1H_1[2
    ],perBankActiveLaneWhenConflict1H_2[2],perBankActiveLaneWhenConflict1H_3[2],perBankActiveLaneWhenConflict1H_4[2],
    perBankActiveLaneWhenConflict1H_5[2],perBankActiveLaneWhenConflict1H_6[2],perBankActiveLaneWhenConflict1H_7[2]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_2 = |_ActiveLaneWhenConflict1H_2_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_3_T_8 = {perBankActiveLaneWhenConflict1H_0[3],perBankActiveLaneWhenConflict1H_1[3
    ],perBankActiveLaneWhenConflict1H_2[3],perBankActiveLaneWhenConflict1H_3[3],perBankActiveLaneWhenConflict1H_4[3],
    perBankActiveLaneWhenConflict1H_5[3],perBankActiveLaneWhenConflict1H_6[3],perBankActiveLaneWhenConflict1H_7[3]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_3 = |_ActiveLaneWhenConflict1H_3_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_4_T_8 = {perBankActiveLaneWhenConflict1H_0[4],perBankActiveLaneWhenConflict1H_1[4
    ],perBankActiveLaneWhenConflict1H_2[4],perBankActiveLaneWhenConflict1H_3[4],perBankActiveLaneWhenConflict1H_4[4],
    perBankActiveLaneWhenConflict1H_5[4],perBankActiveLaneWhenConflict1H_6[4],perBankActiveLaneWhenConflict1H_7[4]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_4 = |_ActiveLaneWhenConflict1H_4_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_5_T_8 = {perBankActiveLaneWhenConflict1H_0[5],perBankActiveLaneWhenConflict1H_1[5
    ],perBankActiveLaneWhenConflict1H_2[5],perBankActiveLaneWhenConflict1H_3[5],perBankActiveLaneWhenConflict1H_4[5],
    perBankActiveLaneWhenConflict1H_5[5],perBankActiveLaneWhenConflict1H_6[5],perBankActiveLaneWhenConflict1H_7[5]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_5 = |_ActiveLaneWhenConflict1H_5_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_6_T_8 = {perBankActiveLaneWhenConflict1H_0[6],perBankActiveLaneWhenConflict1H_1[6
    ],perBankActiveLaneWhenConflict1H_2[6],perBankActiveLaneWhenConflict1H_3[6],perBankActiveLaneWhenConflict1H_4[6],
    perBankActiveLaneWhenConflict1H_5[6],perBankActiveLaneWhenConflict1H_6[6],perBankActiveLaneWhenConflict1H_7[6]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_6 = |_ActiveLaneWhenConflict1H_6_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ActiveLaneWhenConflict1H_7_T_8 = {perBankActiveLaneWhenConflict1H_0[7],perBankActiveLaneWhenConflict1H_1[7
    ],perBankActiveLaneWhenConflict1H_2[7],perBankActiveLaneWhenConflict1H_3[7],perBankActiveLaneWhenConflict1H_4[7],
    perBankActiveLaneWhenConflict1H_5[7],perBankActiveLaneWhenConflict1H_6[7],perBankActiveLaneWhenConflict1H_7[7]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_7 = |_ActiveLaneWhenConflict1H_7_T_8; // @[BankConflictArbiter.scala 156:83]
  wire [7:0] _ReserveLaneWhenConflict1H_T = {ActiveLaneWhenConflict1H_0,ActiveLaneWhenConflict1H_1,
    ActiveLaneWhenConflict1H_2,ActiveLaneWhenConflict1H_3,ActiveLaneWhenConflict1H_4,ActiveLaneWhenConflict1H_5,
    ActiveLaneWhenConflict1H_6,ActiveLaneWhenConflict1H_7}; // @[Cat.scala 31:58]
  wire [7:0] _ReserveLaneWhenConflict1H_T_1 = ~_ReserveLaneWhenConflict1H_T; // @[BankConflictArbiter.scala 157:45]
  wire [7:0] _ReserveLaneWhenConflict1H_T_2 = {perLaneConflictReq_0_activeMask,perLaneConflictReq_1_activeMask,
    perLaneConflictReq_2_activeMask,perLaneConflictReq_3_activeMask,perLaneConflictReq_4_activeMask,
    perLaneConflictReq_5_activeMask,perLaneConflictReq_6_activeMask,perLaneConflictReq_7_activeMask}; // @[Cat.scala 31:58]
  wire [7:0] _ReserveLaneWhenConflict1H_T_3 = _ReserveLaneWhenConflict1H_T_1 & _ReserveLaneWhenConflict1H_T_2; // @[BankConflictArbiter.scala 157:86]
  wire  ReserveLaneWhenConflict1H_7 = _ReserveLaneWhenConflict1H_T_3[0]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_6 = _ReserveLaneWhenConflict1H_T_3[1]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_5 = _ReserveLaneWhenConflict1H_T_3[2]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_4 = _ReserveLaneWhenConflict1H_T_3[3]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_3 = _ReserveLaneWhenConflict1H_T_3[4]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_2 = _ReserveLaneWhenConflict1H_T_3[5]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_1 = _ReserveLaneWhenConflict1H_T_3[6]; // @[BankConflictArbiter.scala 157:109]
  wire  ReserveLaneWhenConflict1H_0 = _ReserveLaneWhenConflict1H_T_3[7]; // @[BankConflictArbiter.scala 157:109]
  wire [3:0] perLaneConflictReq_0_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_0_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_0_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_1_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_1_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_1_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_2_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_2_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_2_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_3_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_3_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_3_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_4_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_4_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_4_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_5_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_5_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_5_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_6_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_6_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_6_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] perLaneConflictReq_7_AddrBundle_wordOffset1H = bankConflict_reg ?
    perLaneConflictReq_reg_7_AddrBundle_wordOffset1H : io_coreReqArb_perLaneAddr_7_wordOffset1H; // @[BankConflictArbiter.scala 159:28]
  wire [3:0] _T_145 = perBankActiveLaneWhenConflict1H_0[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_146 = perBankActiveLaneWhenConflict1H_0[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_147 = perBankActiveLaneWhenConflict1H_0[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_148 = perBankActiveLaneWhenConflict1H_0[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_149 = perBankActiveLaneWhenConflict1H_0[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_150 = perBankActiveLaneWhenConflict1H_0[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_151 = perBankActiveLaneWhenConflict1H_0[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_152 = perBankActiveLaneWhenConflict1H_0[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_153 = _T_145 | _T_146; // @[Mux.scala 27:73]
  wire [3:0] _T_154 = _T_153 | _T_147; // @[Mux.scala 27:73]
  wire [3:0] _T_155 = _T_154 | _T_148; // @[Mux.scala 27:73]
  wire [3:0] _T_156 = _T_155 | _T_149; // @[Mux.scala 27:73]
  wire [3:0] _T_157 = _T_156 | _T_150; // @[Mux.scala 27:73]
  wire [3:0] _T_158 = _T_157 | _T_151; // @[Mux.scala 27:73]
  wire [3:0] _T_168 = perBankActiveLaneWhenConflict1H_1[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_169 = perBankActiveLaneWhenConflict1H_1[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_170 = perBankActiveLaneWhenConflict1H_1[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_171 = perBankActiveLaneWhenConflict1H_1[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_172 = perBankActiveLaneWhenConflict1H_1[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_173 = perBankActiveLaneWhenConflict1H_1[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_174 = perBankActiveLaneWhenConflict1H_1[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_175 = perBankActiveLaneWhenConflict1H_1[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_176 = _T_168 | _T_169; // @[Mux.scala 27:73]
  wire [3:0] _T_177 = _T_176 | _T_170; // @[Mux.scala 27:73]
  wire [3:0] _T_178 = _T_177 | _T_171; // @[Mux.scala 27:73]
  wire [3:0] _T_179 = _T_178 | _T_172; // @[Mux.scala 27:73]
  wire [3:0] _T_180 = _T_179 | _T_173; // @[Mux.scala 27:73]
  wire [3:0] _T_181 = _T_180 | _T_174; // @[Mux.scala 27:73]
  wire [3:0] _T_191 = perBankActiveLaneWhenConflict1H_2[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_192 = perBankActiveLaneWhenConflict1H_2[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_193 = perBankActiveLaneWhenConflict1H_2[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_194 = perBankActiveLaneWhenConflict1H_2[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_195 = perBankActiveLaneWhenConflict1H_2[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_196 = perBankActiveLaneWhenConflict1H_2[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_197 = perBankActiveLaneWhenConflict1H_2[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_198 = perBankActiveLaneWhenConflict1H_2[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_199 = _T_191 | _T_192; // @[Mux.scala 27:73]
  wire [3:0] _T_200 = _T_199 | _T_193; // @[Mux.scala 27:73]
  wire [3:0] _T_201 = _T_200 | _T_194; // @[Mux.scala 27:73]
  wire [3:0] _T_202 = _T_201 | _T_195; // @[Mux.scala 27:73]
  wire [3:0] _T_203 = _T_202 | _T_196; // @[Mux.scala 27:73]
  wire [3:0] _T_204 = _T_203 | _T_197; // @[Mux.scala 27:73]
  wire [3:0] _T_214 = perBankActiveLaneWhenConflict1H_3[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_215 = perBankActiveLaneWhenConflict1H_3[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_216 = perBankActiveLaneWhenConflict1H_3[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_217 = perBankActiveLaneWhenConflict1H_3[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_218 = perBankActiveLaneWhenConflict1H_3[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_219 = perBankActiveLaneWhenConflict1H_3[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_220 = perBankActiveLaneWhenConflict1H_3[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_221 = perBankActiveLaneWhenConflict1H_3[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_222 = _T_214 | _T_215; // @[Mux.scala 27:73]
  wire [3:0] _T_223 = _T_222 | _T_216; // @[Mux.scala 27:73]
  wire [3:0] _T_224 = _T_223 | _T_217; // @[Mux.scala 27:73]
  wire [3:0] _T_225 = _T_224 | _T_218; // @[Mux.scala 27:73]
  wire [3:0] _T_226 = _T_225 | _T_219; // @[Mux.scala 27:73]
  wire [3:0] _T_227 = _T_226 | _T_220; // @[Mux.scala 27:73]
  wire [3:0] _T_237 = perBankActiveLaneWhenConflict1H_4[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_238 = perBankActiveLaneWhenConflict1H_4[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_239 = perBankActiveLaneWhenConflict1H_4[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_240 = perBankActiveLaneWhenConflict1H_4[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_241 = perBankActiveLaneWhenConflict1H_4[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_242 = perBankActiveLaneWhenConflict1H_4[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_243 = perBankActiveLaneWhenConflict1H_4[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_244 = perBankActiveLaneWhenConflict1H_4[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_245 = _T_237 | _T_238; // @[Mux.scala 27:73]
  wire [3:0] _T_246 = _T_245 | _T_239; // @[Mux.scala 27:73]
  wire [3:0] _T_247 = _T_246 | _T_240; // @[Mux.scala 27:73]
  wire [3:0] _T_248 = _T_247 | _T_241; // @[Mux.scala 27:73]
  wire [3:0] _T_249 = _T_248 | _T_242; // @[Mux.scala 27:73]
  wire [3:0] _T_250 = _T_249 | _T_243; // @[Mux.scala 27:73]
  wire [3:0] _T_260 = perBankActiveLaneWhenConflict1H_5[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_261 = perBankActiveLaneWhenConflict1H_5[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_262 = perBankActiveLaneWhenConflict1H_5[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_263 = perBankActiveLaneWhenConflict1H_5[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_264 = perBankActiveLaneWhenConflict1H_5[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_265 = perBankActiveLaneWhenConflict1H_5[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_266 = perBankActiveLaneWhenConflict1H_5[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_267 = perBankActiveLaneWhenConflict1H_5[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_268 = _T_260 | _T_261; // @[Mux.scala 27:73]
  wire [3:0] _T_269 = _T_268 | _T_262; // @[Mux.scala 27:73]
  wire [3:0] _T_270 = _T_269 | _T_263; // @[Mux.scala 27:73]
  wire [3:0] _T_271 = _T_270 | _T_264; // @[Mux.scala 27:73]
  wire [3:0] _T_272 = _T_271 | _T_265; // @[Mux.scala 27:73]
  wire [3:0] _T_273 = _T_272 | _T_266; // @[Mux.scala 27:73]
  wire [3:0] _T_283 = perBankActiveLaneWhenConflict1H_6[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_284 = perBankActiveLaneWhenConflict1H_6[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_285 = perBankActiveLaneWhenConflict1H_6[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_286 = perBankActiveLaneWhenConflict1H_6[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_287 = perBankActiveLaneWhenConflict1H_6[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_288 = perBankActiveLaneWhenConflict1H_6[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_289 = perBankActiveLaneWhenConflict1H_6[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_290 = perBankActiveLaneWhenConflict1H_6[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_291 = _T_283 | _T_284; // @[Mux.scala 27:73]
  wire [3:0] _T_292 = _T_291 | _T_285; // @[Mux.scala 27:73]
  wire [3:0] _T_293 = _T_292 | _T_286; // @[Mux.scala 27:73]
  wire [3:0] _T_294 = _T_293 | _T_287; // @[Mux.scala 27:73]
  wire [3:0] _T_295 = _T_294 | _T_288; // @[Mux.scala 27:73]
  wire [3:0] _T_296 = _T_295 | _T_289; // @[Mux.scala 27:73]
  wire [3:0] _T_306 = perBankActiveLaneWhenConflict1H_7[0] ? perLaneConflictReq_0_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_307 = perBankActiveLaneWhenConflict1H_7[1] ? perLaneConflictReq_1_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_308 = perBankActiveLaneWhenConflict1H_7[2] ? perLaneConflictReq_2_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_309 = perBankActiveLaneWhenConflict1H_7[3] ? perLaneConflictReq_3_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_310 = perBankActiveLaneWhenConflict1H_7[4] ? perLaneConflictReq_4_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_311 = perBankActiveLaneWhenConflict1H_7[5] ? perLaneConflictReq_5_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_312 = perBankActiveLaneWhenConflict1H_7[6] ? perLaneConflictReq_6_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_313 = perBankActiveLaneWhenConflict1H_7[7] ? perLaneConflictReq_7_AddrBundle_wordOffset1H : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_314 = _T_306 | _T_307; // @[Mux.scala 27:73]
  wire [3:0] _T_315 = _T_314 | _T_308; // @[Mux.scala 27:73]
  wire [3:0] _T_316 = _T_315 | _T_309; // @[Mux.scala 27:73]
  wire [3:0] _T_317 = _T_316 | _T_310; // @[Mux.scala 27:73]
  wire [3:0] _T_318 = _T_317 | _T_311; // @[Mux.scala 27:73]
  wire [3:0] _T_319 = _T_318 | _T_312; // @[Mux.scala 27:73]
  assign io_dataCrsbarSel1H_0 = isWrite ? perBankActiveLaneWhenConflict1H_0 : bankIdxMasked_0; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_1 = isWrite ? perBankActiveLaneWhenConflict1H_1 : bankIdxMasked_1; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_2 = isWrite ? perBankActiveLaneWhenConflict1H_2 : bankIdxMasked_2; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_3 = isWrite ? perBankActiveLaneWhenConflict1H_3 : bankIdxMasked_3; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_4 = isWrite ? perBankActiveLaneWhenConflict1H_4 : bankIdxMasked_4; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_5 = isWrite ? perBankActiveLaneWhenConflict1H_5 : bankIdxMasked_5; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_6 = isWrite ? perBankActiveLaneWhenConflict1H_6 : bankIdxMasked_6; // @[BankConflictArbiter.scala 174:28]
  assign io_dataCrsbarSel1H_7 = isWrite ? perBankActiveLaneWhenConflict1H_7 : bankIdxMasked_7; // @[BankConflictArbiter.scala 174:28]
  assign io_addrCrsbarOut_0_wordOffset1H = _T_158 | _T_152; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_1_wordOffset1H = _T_181 | _T_175; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_2_wordOffset1H = _T_204 | _T_198; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_3_wordOffset1H = _T_227 | _T_221; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_4_wordOffset1H = _T_250 | _T_244; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_5_wordOffset1H = _T_273 | _T_267; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_6_wordOffset1H = _T_296 | _T_290; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_7_wordOffset1H = _T_319 | _T_313; // @[Mux.scala 27:73]
  assign io_dataArrayEn_0 = |perBankActiveLaneWhenConflict1H_0; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_1 = |perBankActiveLaneWhenConflict1H_1; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_2 = |perBankActiveLaneWhenConflict1H_2; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_3 = |perBankActiveLaneWhenConflict1H_3; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_4 = |perBankActiveLaneWhenConflict1H_4; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_5 = |perBankActiveLaneWhenConflict1H_5; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_6 = |perBankActiveLaneWhenConflict1H_6; // @[BankConflictArbiter.scala 177:59]
  assign io_dataArrayEn_7 = |perBankActiveLaneWhenConflict1H_7; // @[BankConflictArbiter.scala 177:59]
  assign io_activeLane_0 = |_ActiveLaneWhenConflict1H_0_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_1 = |_ActiveLaneWhenConflict1H_1_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_2 = |_ActiveLaneWhenConflict1H_2_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_3 = |_ActiveLaneWhenConflict1H_3_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_4 = |_ActiveLaneWhenConflict1H_4_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_5 = |_ActiveLaneWhenConflict1H_5_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_6 = |_ActiveLaneWhenConflict1H_6_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_activeLane_7 = |_ActiveLaneWhenConflict1H_7_T_8; // @[BankConflictArbiter.scala 156:83]
  assign io_bankConflict = |_bankConflict_T & (io_coreReqArb_enable | bankConflict_reg); // @[BankConflictArbiter.scala 148:47]
  always @(posedge clock) begin
    if (reset) begin // @[BankConflictArbiter.scala 105:33]
      bankConflict_reg <= 1'h0; // @[BankConflictArbiter.scala 105:33]
    end else begin
      bankConflict_reg <= bankConflict; // @[BankConflictArbiter.scala 105:33]
    end
    if (bankConflict) begin // @[BankConflictArbiter.scala 167:21]
      conflictReqIsW_reg <= io_coreReqArb_isWrite; // @[BankConflictArbiter.scala 167:41]
    end
    perLaneConflictReq_reg_0_activeMask <= _ReserveLaneWhenConflict1H_T_3[7]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_0) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_0_bankIdx <= io_coreReqArb_perLaneAddr_0_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_0) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_0_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_0_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_1_activeMask <= _ReserveLaneWhenConflict1H_T_3[6]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_1) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_1_bankIdx <= io_coreReqArb_perLaneAddr_1_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_1) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_1_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_1_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_2_activeMask <= _ReserveLaneWhenConflict1H_T_3[5]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_2) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_2_bankIdx <= io_coreReqArb_perLaneAddr_2_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_2) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_2_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_2_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_3_activeMask <= _ReserveLaneWhenConflict1H_T_3[4]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_3) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_3_bankIdx <= io_coreReqArb_perLaneAddr_3_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_3) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_3_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_3_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_4_activeMask <= _ReserveLaneWhenConflict1H_T_3[3]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_4) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_4_bankIdx <= io_coreReqArb_perLaneAddr_4_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_4) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_4_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_4_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_5_activeMask <= _ReserveLaneWhenConflict1H_T_3[2]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_5) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_5_bankIdx <= io_coreReqArb_perLaneAddr_5_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_5) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_5_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_5_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_6_activeMask <= _ReserveLaneWhenConflict1H_T_3[1]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_6) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_6_bankIdx <= io_coreReqArb_perLaneAddr_6_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_6) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_6_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_6_wordOffset1H;
      end
    end
    perLaneConflictReq_reg_7_activeMask <= _ReserveLaneWhenConflict1H_T_3[0]; // @[BankConflictArbiter.scala 157:109]
    if (ReserveLaneWhenConflict1H_7) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_7_bankIdx <= io_coreReqArb_perLaneAddr_7_blockOffset;
      end
    end
    if (ReserveLaneWhenConflict1H_7) begin // @[BankConflictArbiter.scala 162:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 159:28]
        perLaneConflictReq_reg_7_AddrBundle_wordOffset1H <= io_coreReqArb_perLaneAddr_7_wordOffset1H;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bankConflict_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  conflictReqIsW_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  perLaneConflictReq_reg_0_activeMask = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  perLaneConflictReq_reg_0_bankIdx = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  perLaneConflictReq_reg_0_AddrBundle_wordOffset1H = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  perLaneConflictReq_reg_1_activeMask = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  perLaneConflictReq_reg_1_bankIdx = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  perLaneConflictReq_reg_1_AddrBundle_wordOffset1H = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  perLaneConflictReq_reg_2_activeMask = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  perLaneConflictReq_reg_2_bankIdx = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  perLaneConflictReq_reg_2_AddrBundle_wordOffset1H = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  perLaneConflictReq_reg_3_activeMask = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  perLaneConflictReq_reg_3_bankIdx = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  perLaneConflictReq_reg_3_AddrBundle_wordOffset1H = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  perLaneConflictReq_reg_4_activeMask = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  perLaneConflictReq_reg_4_bankIdx = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  perLaneConflictReq_reg_4_AddrBundle_wordOffset1H = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  perLaneConflictReq_reg_5_activeMask = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  perLaneConflictReq_reg_5_bankIdx = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  perLaneConflictReq_reg_5_AddrBundle_wordOffset1H = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  perLaneConflictReq_reg_6_activeMask = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  perLaneConflictReq_reg_6_bankIdx = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  perLaneConflictReq_reg_6_AddrBundle_wordOffset1H = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  perLaneConflictReq_reg_7_activeMask = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  perLaneConflictReq_reg_7_bankIdx = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  perLaneConflictReq_reg_7_AddrBundle_wordOffset1H = _RAND_25[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MSHR_1(
  input         clock,
  input         reset,
  output        io_missReq_ready,
  input         io_missReq_valid,
  input  [26:0] io_missReq_bits_blockAddr,
  input  [1:0]  io_missReq_bits_instrId,
  input  [64:0] io_missReq_bits_targetInfo,
  output        io_missRspIn_ready,
  input         io_missRspIn_valid,
  input  [26:0] io_missRspIn_bits_blockAddr,
  input         io_missRspOut_ready,
  output        io_missRspOut_valid,
  output [64:0] io_missRspOut_bits_targetInfo,
  output [26:0] io_missRspOut_bits_blockAddr,
  output [1:0]  io_missRspOut_bits_instrId,
  input         io_miss2mem_ready,
  output        io_miss2mem_valid,
  output [26:0] io_miss2mem_bits_blockAddr,
  output [1:0]  io_miss2mem_bits_instrId
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [95:0] _RAND_20;
  reg [95:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [95:0] _RAND_24;
  reg [95:0] _RAND_25;
  reg [95:0] _RAND_26;
  reg [95:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [95:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [95:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] subentryStatus_io_valid_list; // @[DCacheMSHR.scala 77:30]
  wire  subentryStatus_io_full; // @[DCacheMSHR.scala 77:30]
  wire [1:0] subentryStatus_io_next; // @[DCacheMSHR.scala 77:30]
  wire [2:0] subentryStatus_io_used; // @[DCacheMSHR.scala 77:30]
  wire [3:0] entryStatus_io_valid_list; // @[DCacheMSHR.scala 84:27]
  wire  entryStatus_io_full; // @[DCacheMSHR.scala 84:27]
  wire [1:0] entryStatus_io_next; // @[DCacheMSHR.scala 84:27]
  wire [2:0] entryStatus_io_used; // @[DCacheMSHR.scala 84:27]
  wire [3:0] hasSendStatus_io_valid_list; // @[DCacheMSHR.scala 156:29]
  wire  hasSendStatus_io_full; // @[DCacheMSHR.scala 156:29]
  wire [1:0] hasSendStatus_io_next; // @[DCacheMSHR.scala 156:29]
  wire [2:0] hasSendStatus_io_used; // @[DCacheMSHR.scala 156:29]
  reg [26:0] blockAddr_Access_0; // @[DCacheMSHR.scala 51:33]
  reg [26:0] blockAddr_Access_1; // @[DCacheMSHR.scala 51:33]
  reg [26:0] blockAddr_Access_2; // @[DCacheMSHR.scala 51:33]
  reg [26:0] blockAddr_Access_3; // @[DCacheMSHR.scala 51:33]
  reg [1:0] instrId_Access_0_0; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_0_1; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_0_2; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_0_3; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_1_0; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_1_1; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_1_2; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_1_3; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_2_0; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_2_1; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_2_2; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_2_3; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_3_0; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_3_1; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_3_2; // @[DCacheMSHR.scala 52:31]
  reg [1:0] instrId_Access_3_3; // @[DCacheMSHR.scala 52:31]
  reg [64:0] targetInfo_Accesss_0_0; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_0_1; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_0_2; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_0_3; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_1_0; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_1_1; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_1_2; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_1_3; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_2_0; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_2_1; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_2_2; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_2_3; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_3_0; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_3_1; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_3_2; // @[DCacheMSHR.scala 53:35]
  reg [64:0] targetInfo_Accesss_3_3; // @[DCacheMSHR.scala 53:35]
  reg  subentry_valid_0_0; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_0_1; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_0_2; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_0_3; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_1_0; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_1_1; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_1_2; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_1_3; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_2_0; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_2_1; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_2_2; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_2_3; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_3_0; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_3_1; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_3_2; // @[DCacheMSHR.scala 75:31]
  reg  subentry_valid_3_3; // @[DCacheMSHR.scala 75:31]
  wire  _entryMatchMissRsp_T = blockAddr_Access_0 == io_missRspIn_bits_blockAddr; // @[DCacheMSHR.scala 87:58]
  wire  _entryMatchMissRsp_T_1 = blockAddr_Access_1 == io_missRspIn_bits_blockAddr; // @[DCacheMSHR.scala 87:58]
  wire  _entryMatchMissRsp_T_2 = blockAddr_Access_2 == io_missRspIn_bits_blockAddr; // @[DCacheMSHR.scala 87:58]
  wire  _entryMatchMissRsp_T_3 = blockAddr_Access_3 == io_missRspIn_bits_blockAddr; // @[DCacheMSHR.scala 87:58]
  wire [3:0] _entryMatchMissRsp_T_4 = {_entryMatchMissRsp_T,_entryMatchMissRsp_T_1,_entryMatchMissRsp_T_2,
    _entryMatchMissRsp_T_3}; // @[Cat.scala 31:58]
  wire [3:0] _entryMatchMissRsp_T_13 = {_entryMatchMissRsp_T_4[0],_entryMatchMissRsp_T_4[1],_entryMatchMissRsp_T_4[2],
    _entryMatchMissRsp_T_4[3]}; // @[Cat.scala 31:58]
  wire [3:0] _entry_valid_T = {subentry_valid_0_0,subentry_valid_0_1,subentry_valid_0_2,subentry_valid_0_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_1 = |_entry_valid_T; // @[DCacheMSHR.scala 83:59]
  wire [3:0] _entry_valid_T_2 = {subentry_valid_1_0,subentry_valid_1_1,subentry_valid_1_2,subentry_valid_1_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_3 = |_entry_valid_T_2; // @[DCacheMSHR.scala 83:59]
  wire [3:0] _entry_valid_T_4 = {subentry_valid_2_0,subentry_valid_2_1,subentry_valid_2_2,subentry_valid_2_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_5 = |_entry_valid_T_4; // @[DCacheMSHR.scala 83:59]
  wire [3:0] _entry_valid_T_6 = {subentry_valid_3_0,subentry_valid_3_1,subentry_valid_3_2,subentry_valid_3_3}; // @[Cat.scala 31:58]
  wire  _entry_valid_T_7 = |_entry_valid_T_6; // @[DCacheMSHR.scala 83:59]
  wire [3:0] _entry_valid_T_8 = {_entry_valid_T_1,_entry_valid_T_3,_entry_valid_T_5,_entry_valid_T_7}; // @[Cat.scala 31:58]
  wire [1:0] _entry_valid_T_12 = {_entry_valid_T_8[0],_entry_valid_T_8[1]}; // @[Cat.scala 31:58]
  wire [1:0] _entry_valid_T_16 = {_entry_valid_T_8[2],_entry_valid_T_8[3]}; // @[Cat.scala 31:58]
  wire [3:0] entry_valid = {_entry_valid_T_8[0],_entry_valid_T_8[1],_entry_valid_T_8[2],_entry_valid_T_8[3]}; // @[Cat.scala 31:58]
  wire [3:0] entryMatchMissRsp = _entryMatchMissRsp_T_13 & entry_valid; // @[DCacheMSHR.scala 87:92]
  wire [1:0] subentry_selected_hi = entryMatchMissRsp[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] subentry_selected_lo = entryMatchMissRsp[1:0]; // @[OneHot.scala 31:18]
  wire  _subentry_selected_T = |subentry_selected_hi; // @[OneHot.scala 32:14]
  wire [1:0] _subentry_selected_T_1 = subentry_selected_hi | subentry_selected_lo; // @[OneHot.scala 32:28]
  wire [1:0] _subentry_selected_T_3 = {_subentry_selected_T,_subentry_selected_T_1[1]}; // @[Cat.scala 31:58]
  wire  _GEN_1 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_2 : subentry_valid_0_2; // @[Cat.scala 31:{58,58}]
  wire  _GEN_2 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_2 : _GEN_1; // @[Cat.scala 31:{58,58}]
  wire  _GEN_3 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_2 : _GEN_2; // @[Cat.scala 31:{58,58}]
  wire  _GEN_5 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_3 : subentry_valid_0_3; // @[Cat.scala 31:{58,58}]
  wire  _GEN_6 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_3 : _GEN_5; // @[Cat.scala 31:{58,58}]
  wire  _GEN_7 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_3 : _GEN_6; // @[Cat.scala 31:{58,58}]
  wire  _GEN_9 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_0 : subentry_valid_0_0; // @[Cat.scala 31:{58,58}]
  wire  _GEN_10 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_0 : _GEN_9; // @[Cat.scala 31:{58,58}]
  wire  _GEN_11 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_0 : _GEN_10; // @[Cat.scala 31:{58,58}]
  wire  _GEN_13 = 2'h1 == _subentry_selected_T_3 ? subentry_valid_1_1 : subentry_valid_0_1; // @[Cat.scala 31:{58,58}]
  wire  _GEN_14 = 2'h2 == _subentry_selected_T_3 ? subentry_valid_2_1 : _GEN_13; // @[Cat.scala 31:{58,58}]
  wire  _GEN_15 = 2'h3 == _subentry_selected_T_3 ? subentry_valid_3_1 : _GEN_14; // @[Cat.scala 31:{58,58}]
  wire [3:0] _subentryStatus_io_valid_list_T = {_GEN_11,_GEN_15,_GEN_3,_GEN_7}; // @[Cat.scala 31:58]
  wire [1:0] _subentryStatus_io_valid_list_T_4 = {_subentryStatus_io_valid_list_T[0],_subentryStatus_io_valid_list_T[1]}
    ; // @[Cat.scala 31:58]
  wire [1:0] _subentryStatus_io_valid_list_T_8 = {_subentryStatus_io_valid_list_T[2],_subentryStatus_io_valid_list_T[3]}
    ; // @[Cat.scala 31:58]
  wire [1:0] _subentry_next2cancel_T_4 = _GEN_3 ? 2'h2 : 2'h3; // @[DCacheMSHR.scala 80:55]
  wire [1:0] _subentry_next2cancel_T_5 = _GEN_15 ? 2'h1 : _subentry_next2cancel_T_4; // @[DCacheMSHR.scala 80:55]
  wire [1:0] subentry_next2cancel = _GEN_11 ? 2'h0 : _subentry_next2cancel_T_5; // @[DCacheMSHR.scala 80:55]
  wire [1:0] _T_4 = entryMatchMissRsp[0] + entryMatchMissRsp[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _T_6 = entryMatchMissRsp[2] + entryMatchMissRsp[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _T_8 = _T_4 + _T_6; // @[Bitwise.scala 48:55]
  wire  _T_12 = ~reset; // @[DCacheMSHR.scala 88:9]
  wire  _entryMatchMissReq_T = blockAddr_Access_0 == io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 89:58]
  wire  _entryMatchMissReq_T_1 = blockAddr_Access_1 == io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 89:58]
  wire  _entryMatchMissReq_T_2 = blockAddr_Access_2 == io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 89:58]
  wire  _entryMatchMissReq_T_3 = blockAddr_Access_3 == io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 89:58]
  wire [3:0] _entryMatchMissReq_T_4 = {_entryMatchMissReq_T,_entryMatchMissReq_T_1,_entryMatchMissReq_T_2,
    _entryMatchMissReq_T_3}; // @[Cat.scala 31:58]
  wire [3:0] _entryMatchMissReq_T_13 = {_entryMatchMissReq_T_4[0],_entryMatchMissReq_T_4[1],_entryMatchMissReq_T_4[2],
    _entryMatchMissReq_T_4[3]}; // @[Cat.scala 31:58]
  wire [3:0] entryMatchMissReq = _entryMatchMissReq_T_13 & entry_valid; // @[DCacheMSHR.scala 89:90]
  wire [1:0] _T_18 = entryMatchMissReq[0] + entryMatchMissReq[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _T_20 = entryMatchMissReq[2] + entryMatchMissReq[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _T_22 = _T_18 + _T_20; // @[Bitwise.scala 48:55]
  wire  secondary_miss = |entryMatchMissReq; // @[DCacheMSHR.scala 92:42]
  wire  primary_miss = ~secondary_miss; // @[DCacheMSHR.scala 93:22]
  reg  missRspBusy; // @[DCacheMSHR.scala 96:28]
  wire  _io_missReq_ready_T_3 = subentryStatus_io_full & secondary_miss; // @[DCacheMSHR.scala 98:29]
  wire  missReq_fire = io_missReq_ready & io_missReq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] real_SRAMAddrUp_hi = entryMatchMissReq[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] real_SRAMAddrUp_lo = entryMatchMissReq[1:0]; // @[OneHot.scala 31:18]
  wire  _real_SRAMAddrUp_T = |real_SRAMAddrUp_hi; // @[OneHot.scala 32:14]
  wire [1:0] _real_SRAMAddrUp_T_1 = real_SRAMAddrUp_hi | real_SRAMAddrUp_lo; // @[OneHot.scala 32:28]
  wire [1:0] _real_SRAMAddrUp_T_3 = {_real_SRAMAddrUp_T,_real_SRAMAddrUp_T_1[1]}; // @[Cat.scala 31:58]
  wire [1:0] real_SRAMAddrUp = secondary_miss ? _real_SRAMAddrUp_T_3 : entryStatus_io_next; // @[DCacheMSHR.scala 103:28]
  wire [1:0] real_SRAMAddrDown = secondary_miss ? subentryStatus_io_next : 2'h0; // @[DCacheMSHR.scala 104:30]
  wire  _T_28 = io_missRspIn_ready & io_missRspIn_valid; // @[Decoupled.scala 50:35]
  wire  _T_42 = subentryStatus_io_used == 3'h1; // @[DCacheMSHR.scala 118:52]
  wire  _GEN_48 = missRspBusy & subentryStatus_io_used == 3'h1 & io_missRspOut_ready ? 1'h0 : missRspBusy; // @[DCacheMSHR.scala 118:83 119:17 96:28]
  wire  _GEN_49 = _T_28 & (subentryStatus_io_used != 3'h1 | ~io_missRspOut_ready) | _GEN_48; // @[DCacheMSHR.scala 116:86 117:17]
  wire  _GEN_252 = 2'h0 == _subentry_selected_T_3; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_253 = 2'h1 == subentry_next2cancel; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_51 = 2'h0 == _subentry_selected_T_3 & 2'h1 == subentry_next2cancel ? targetInfo_Accesss_0_1 :
    targetInfo_Accesss_0_0; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_255 = 2'h2 == subentry_next2cancel; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_52 = 2'h0 == _subentry_selected_T_3 & 2'h2 == subentry_next2cancel ? targetInfo_Accesss_0_2 : _GEN_51
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_257 = 2'h3 == subentry_next2cancel; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_53 = 2'h0 == _subentry_selected_T_3 & 2'h3 == subentry_next2cancel ? targetInfo_Accesss_0_3 : _GEN_52
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_258 = 2'h1 == _subentry_selected_T_3; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_259 = 2'h0 == subentry_next2cancel; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_54 = 2'h1 == _subentry_selected_T_3 & 2'h0 == subentry_next2cancel ? targetInfo_Accesss_1_0 : _GEN_53
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_55 = 2'h1 == _subentry_selected_T_3 & 2'h1 == subentry_next2cancel ? targetInfo_Accesss_1_1 : _GEN_54
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_56 = 2'h1 == _subentry_selected_T_3 & 2'h2 == subentry_next2cancel ? targetInfo_Accesss_1_2 : _GEN_55
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_57 = 2'h1 == _subentry_selected_T_3 & 2'h3 == subentry_next2cancel ? targetInfo_Accesss_1_3 : _GEN_56
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_266 = 2'h2 == _subentry_selected_T_3; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_58 = 2'h2 == _subentry_selected_T_3 & 2'h0 == subentry_next2cancel ? targetInfo_Accesss_2_0 : _GEN_57
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_59 = 2'h2 == _subentry_selected_T_3 & 2'h1 == subentry_next2cancel ? targetInfo_Accesss_2_1 : _GEN_58
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_60 = 2'h2 == _subentry_selected_T_3 & 2'h2 == subentry_next2cancel ? targetInfo_Accesss_2_2 : _GEN_59
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_61 = 2'h2 == _subentry_selected_T_3 & 2'h3 == subentry_next2cancel ? targetInfo_Accesss_2_3 : _GEN_60
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire  _GEN_274 = 2'h3 == _subentry_selected_T_3; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_62 = 2'h3 == _subentry_selected_T_3 & 2'h0 == subentry_next2cancel ? targetInfo_Accesss_3_0 : _GEN_61
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_63 = 2'h3 == _subentry_selected_T_3 & 2'h1 == subentry_next2cancel ? targetInfo_Accesss_3_1 : _GEN_62
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [64:0] _GEN_64 = 2'h3 == _subentry_selected_T_3 & 2'h2 == subentry_next2cancel ? targetInfo_Accesss_3_2 : _GEN_63
    ; // @[DCacheMSHR.scala 123:{33,33}]
  wire [26:0] _GEN_67 = 2'h1 == _subentry_selected_T_3 ? blockAddr_Access_1 : blockAddr_Access_0; // @[DCacheMSHR.scala 124:{32,32}]
  wire [26:0] _GEN_68 = 2'h2 == _subentry_selected_T_3 ? blockAddr_Access_2 : _GEN_67; // @[DCacheMSHR.scala 124:{32,32}]
  wire  _T_45 = 2'h0 == entryStatus_io_next; // @[DCacheMSHR.scala 132:24]
  wire  _T_56 = io_missRspOut_ready & io_missRspOut_valid; // @[Decoupled.scala 50:35]
  wire  _T_57 = _GEN_259 & _T_56; // @[DCacheMSHR.scala 136:53]
  wire  _T_58 = 2'h0 == subentryStatus_io_next; // @[DCacheMSHR.scala 139:35]
  wire  _T_59 = 2'h0 == subentryStatus_io_next & missReq_fire; // @[DCacheMSHR.scala 139:61]
  wire  _GEN_70 = _T_59 & secondary_miss | subentry_valid_0_0; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_71 = _T_57 ? 1'h0 : _GEN_70; // @[DCacheMSHR.scala 137:32 138:43]
  wire  _GEN_72 = _GEN_252 ? _GEN_71 : subentry_valid_0_0; // @[DCacheMSHR.scala 135:61 75:31]
  wire  _GEN_73 = _T_45 & missReq_fire & primary_miss | _GEN_72; // @[DCacheMSHR.scala 133:63 134:41]
  wire  _T_73 = _GEN_253 & _T_56; // @[DCacheMSHR.scala 136:53]
  wire  _T_74 = 2'h1 == subentryStatus_io_next; // @[DCacheMSHR.scala 139:35]
  wire  _T_75 = 2'h1 == subentryStatus_io_next & missReq_fire; // @[DCacheMSHR.scala 139:61]
  wire  _GEN_74 = _T_75 & secondary_miss | subentry_valid_0_1; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _T_89 = _GEN_255 & _T_56; // @[DCacheMSHR.scala 136:53]
  wire  _T_90 = 2'h2 == subentryStatus_io_next; // @[DCacheMSHR.scala 139:35]
  wire  _T_91 = 2'h2 == subentryStatus_io_next & missReq_fire; // @[DCacheMSHR.scala 139:61]
  wire  _GEN_78 = _T_91 & secondary_miss | subentry_valid_0_2; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _T_105 = _GEN_257 & _T_56; // @[DCacheMSHR.scala 136:53]
  wire  _T_106 = 2'h3 == subentryStatus_io_next; // @[DCacheMSHR.scala 139:35]
  wire  _T_107 = 2'h3 == subentryStatus_io_next & missReq_fire; // @[DCacheMSHR.scala 139:61]
  wire  _GEN_82 = _T_107 & secondary_miss | subentry_valid_0_3; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _T_109 = 2'h1 == entryStatus_io_next; // @[DCacheMSHR.scala 132:24]
  wire  _GEN_86 = _T_59 & secondary_miss | subentry_valid_1_0; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_87 = _T_57 ? 1'h0 : _GEN_86; // @[DCacheMSHR.scala 137:32 138:43]
  wire  _GEN_88 = _GEN_258 ? _GEN_87 : subentry_valid_1_0; // @[DCacheMSHR.scala 135:61 75:31]
  wire  _GEN_89 = _T_109 & missReq_fire & primary_miss | _GEN_88; // @[DCacheMSHR.scala 133:63 134:41]
  wire  _GEN_90 = _T_75 & secondary_miss | subentry_valid_1_1; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_94 = _T_91 & secondary_miss | subentry_valid_1_2; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_98 = _T_107 & secondary_miss | subentry_valid_1_3; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _T_173 = 2'h2 == entryStatus_io_next; // @[DCacheMSHR.scala 132:24]
  wire  _GEN_102 = _T_59 & secondary_miss | subentry_valid_2_0; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_103 = _T_57 ? 1'h0 : _GEN_102; // @[DCacheMSHR.scala 137:32 138:43]
  wire  _GEN_104 = _GEN_266 ? _GEN_103 : subentry_valid_2_0; // @[DCacheMSHR.scala 135:61 75:31]
  wire  _GEN_105 = _T_173 & missReq_fire & primary_miss | _GEN_104; // @[DCacheMSHR.scala 133:63 134:41]
  wire  _GEN_106 = _T_75 & secondary_miss | subentry_valid_2_1; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_110 = _T_91 & secondary_miss | subentry_valid_2_2; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_114 = _T_107 & secondary_miss | subentry_valid_2_3; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _T_237 = 2'h3 == entryStatus_io_next; // @[DCacheMSHR.scala 132:24]
  wire  _GEN_118 = _T_59 & secondary_miss | subentry_valid_3_0; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_119 = _T_57 ? 1'h0 : _GEN_118; // @[DCacheMSHR.scala 137:32 138:43]
  wire  _GEN_120 = _GEN_274 ? _GEN_119 : subentry_valid_3_0; // @[DCacheMSHR.scala 135:61 75:31]
  wire  _GEN_121 = _T_237 & missReq_fire & primary_miss | _GEN_120; // @[DCacheMSHR.scala 133:63 134:41]
  wire  _GEN_122 = _T_75 & secondary_miss | subentry_valid_3_1; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_126 = _T_91 & secondary_miss | subentry_valid_3_2; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  wire  _GEN_130 = _T_107 & secondary_miss | subentry_valid_3_3; // @[DCacheMSHR.scala 140:42 141:43 75:31]
  reg  has_send2mem_0; // @[DCacheMSHR.scala 155:29]
  reg  has_send2mem_1; // @[DCacheMSHR.scala 155:29]
  reg  has_send2mem_2; // @[DCacheMSHR.scala 155:29]
  reg  has_send2mem_3; // @[DCacheMSHR.scala 155:29]
  wire [3:0] _hasSendStatus_io_valid_list_T = {has_send2mem_0,has_send2mem_1,has_send2mem_2,has_send2mem_3}; // @[Cat.scala 31:58]
  wire [1:0] _hasSendStatus_io_valid_list_T_4 = {_hasSendStatus_io_valid_list_T[0],_hasSendStatus_io_valid_list_T[1]}; // @[Cat.scala 31:58]
  wire [1:0] _hasSendStatus_io_valid_list_T_8 = {_hasSendStatus_io_valid_list_T[2],_hasSendStatus_io_valid_list_T[3]}; // @[Cat.scala 31:58]
  wire  _GEN_187 = 2'h1 == hasSendStatus_io_next ? has_send2mem_1 : has_send2mem_0; // @[DCacheMSHR.scala 158:{24,24}]
  wire  _GEN_188 = 2'h2 == hasSendStatus_io_next ? has_send2mem_2 : _GEN_187; // @[DCacheMSHR.scala 158:{24,24}]
  wire  _GEN_189 = 2'h3 == hasSendStatus_io_next ? has_send2mem_3 : _GEN_188; // @[DCacheMSHR.scala 158:{24,24}]
  wire [3:0] _io_miss2mem_valid_T_1 = entry_valid >> hasSendStatus_io_next; // @[DCacheMSHR.scala 158:75]
  wire  miss2mem_fire = io_miss2mem_valid & io_miss2mem_ready; // @[DCacheMSHR.scala 159:41]
  wire  _GEN_190 = _T_56 & _T_42 & _GEN_252 ? 1'h0 : has_send2mem_0; // @[DCacheMSHR.scala 164:108 165:25 155:29]
  wire  _GEN_191 = miss2mem_fire & 2'h0 == hasSendStatus_io_next | _GEN_190; // @[DCacheMSHR.scala 162:57 163:25]
  wire  _GEN_192 = _T_56 & _T_42 & _GEN_258 ? 1'h0 : has_send2mem_1; // @[DCacheMSHR.scala 164:108 165:25 155:29]
  wire  _GEN_193 = miss2mem_fire & 2'h1 == hasSendStatus_io_next | _GEN_192; // @[DCacheMSHR.scala 162:57 163:25]
  wire  _GEN_194 = _T_56 & _T_42 & _GEN_266 ? 1'h0 : has_send2mem_2; // @[DCacheMSHR.scala 164:108 165:25 155:29]
  wire  _GEN_195 = miss2mem_fire & 2'h2 == hasSendStatus_io_next | _GEN_194; // @[DCacheMSHR.scala 162:57 163:25]
  wire  _GEN_196 = _T_56 & _T_42 & _GEN_274 ? 1'h0 : has_send2mem_3; // @[DCacheMSHR.scala 164:108 165:25 155:29]
  wire  _GEN_197 = miss2mem_fire & 2'h3 == hasSendStatus_io_next | _GEN_196; // @[DCacheMSHR.scala 162:57 163:25]
  wire [2:0] _GEN_314 = {{1'd0}, hasSendStatus_io_next}; // @[DCacheMSHR.scala 162:31]
  wire [2:0] _GEN_315 = {{1'd0}, _subentry_selected_T_3}; // @[DCacheMSHR.scala 164:76]
  wire  _GEN_198 = _T_56 & _T_42 & 3'h4 == _GEN_315 ? 1'h0 : _GEN_191; // @[DCacheMSHR.scala 164:108 165:25]
  wire  _GEN_199 = miss2mem_fire & 3'h4 == _GEN_314 | _GEN_198; // @[DCacheMSHR.scala 162:57 163:25]
  wire  _rInstrId_T = missRspBusy | io_missRspIn_valid; // @[DCacheMSHR.scala 168:46]
  wire [1:0] _rInstrId_T_5 = missRspBusy | io_missRspIn_valid ? _subentry_selected_T_3 : hasSendStatus_io_next; // @[DCacheMSHR.scala 168:33]
  wire [1:0] _rInstrId_T_7 = _rInstrId_T ? subentry_next2cancel : 2'h0; // @[DCacheMSHR.scala 169:60]
  wire [1:0] _GEN_201 = 2'h0 == _rInstrId_T_5 & 2'h1 == _rInstrId_T_7 ? instrId_Access_0_1 : instrId_Access_0_0; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_202 = 2'h0 == _rInstrId_T_5 & 2'h2 == _rInstrId_T_7 ? instrId_Access_0_2 : _GEN_201; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_203 = 2'h0 == _rInstrId_T_5 & 2'h3 == _rInstrId_T_7 ? instrId_Access_0_3 : _GEN_202; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_204 = 2'h1 == _rInstrId_T_5 & 2'h0 == _rInstrId_T_7 ? instrId_Access_1_0 : _GEN_203; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_205 = 2'h1 == _rInstrId_T_5 & 2'h1 == _rInstrId_T_7 ? instrId_Access_1_1 : _GEN_204; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_206 = 2'h1 == _rInstrId_T_5 & 2'h2 == _rInstrId_T_7 ? instrId_Access_1_2 : _GEN_205; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_207 = 2'h1 == _rInstrId_T_5 & 2'h3 == _rInstrId_T_7 ? instrId_Access_1_3 : _GEN_206; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_208 = 2'h2 == _rInstrId_T_5 & 2'h0 == _rInstrId_T_7 ? instrId_Access_2_0 : _GEN_207; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_209 = 2'h2 == _rInstrId_T_5 & 2'h1 == _rInstrId_T_7 ? instrId_Access_2_1 : _GEN_208; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_210 = 2'h2 == _rInstrId_T_5 & 2'h2 == _rInstrId_T_7 ? instrId_Access_2_2 : _GEN_209; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_211 = 2'h2 == _rInstrId_T_5 & 2'h3 == _rInstrId_T_7 ? instrId_Access_2_3 : _GEN_210; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_212 = 2'h3 == _rInstrId_T_5 & 2'h0 == _rInstrId_T_7 ? instrId_Access_3_0 : _GEN_211; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_213 = 2'h3 == _rInstrId_T_5 & 2'h1 == _rInstrId_T_7 ? instrId_Access_3_1 : _GEN_212; // @[DCacheMSHR.scala 168:{12,12}]
  wire [1:0] _GEN_214 = 2'h3 == _rInstrId_T_5 & 2'h2 == _rInstrId_T_7 ? instrId_Access_3_2 : _GEN_213; // @[DCacheMSHR.scala 168:{12,12}]
  wire [26:0] _GEN_217 = 2'h1 == hasSendStatus_io_next ? blockAddr_Access_1 : blockAddr_Access_0; // @[DCacheMSHR.scala 170:{30,30}]
  wire [26:0] _GEN_218 = 2'h2 == hasSendStatus_io_next ? blockAddr_Access_2 : _GEN_217; // @[DCacheMSHR.scala 170:{30,30}]
  getEntryStatus subentryStatus ( // @[DCacheMSHR.scala 77:30]
    .io_valid_list(subentryStatus_io_valid_list),
    .io_full(subentryStatus_io_full),
    .io_next(subentryStatus_io_next),
    .io_used(subentryStatus_io_used)
  );
  getEntryStatus entryStatus ( // @[DCacheMSHR.scala 84:27]
    .io_valid_list(entryStatus_io_valid_list),
    .io_full(entryStatus_io_full),
    .io_next(entryStatus_io_next),
    .io_used(entryStatus_io_used)
  );
  getEntryStatus hasSendStatus ( // @[DCacheMSHR.scala 156:29]
    .io_valid_list(hasSendStatus_io_valid_list),
    .io_full(hasSendStatus_io_full),
    .io_next(hasSendStatus_io_next),
    .io_used(hasSendStatus_io_used)
  );
  assign io_missReq_ready = ~((entryStatus_io_full | missRspBusy | io_missRspIn_valid) & primary_miss |
    _io_missReq_ready_T_3); // @[DCacheMSHR.scala 97:23]
  assign io_missRspIn_ready = ~missRspBusy & io_missRspOut_ready; // @[DCacheMSHR.scala 121:38]
  assign io_missRspOut_valid = io_missRspIn_valid | missRspBusy; // @[DCacheMSHR.scala 127:45]
  assign io_missRspOut_bits_targetInfo = 2'h3 == _subentry_selected_T_3 & 2'h3 == subentry_next2cancel ?
    targetInfo_Accesss_3_3 : _GEN_64; // @[DCacheMSHR.scala 123:{33,33}]
  assign io_missRspOut_bits_blockAddr = 2'h3 == _subentry_selected_T_3 ? blockAddr_Access_3 : _GEN_68; // @[DCacheMSHR.scala 124:{32,32}]
  assign io_missRspOut_bits_instrId = 2'h3 == _rInstrId_T_5 & 2'h3 == _rInstrId_T_7 ? instrId_Access_3_3 : _GEN_214; // @[DCacheMSHR.scala 168:{12,12}]
  assign io_miss2mem_valid = ~_GEN_189 & _io_miss2mem_valid_T_1[0]; // @[DCacheMSHR.scala 158:61]
  assign io_miss2mem_bits_blockAddr = 2'h3 == hasSendStatus_io_next ? blockAddr_Access_3 : _GEN_218; // @[DCacheMSHR.scala 170:{30,30}]
  assign io_miss2mem_bits_instrId = 2'h3 == _rInstrId_T_5 & 2'h3 == _rInstrId_T_7 ? instrId_Access_3_3 : _GEN_214; // @[DCacheMSHR.scala 168:{12,12}]
  assign subentryStatus_io_valid_list = {_subentryStatus_io_valid_list_T_4,_subentryStatus_io_valid_list_T_8}; // @[Cat.scala 31:58]
  assign entryStatus_io_valid_list = {_entry_valid_T_12,_entry_valid_T_16}; // @[Cat.scala 31:58]
  assign hasSendStatus_io_valid_list = {_hasSendStatus_io_valid_list_T_4,_hasSendStatus_io_valid_list_T_8}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[DCacheMSHR.scala 51:33]
      blockAddr_Access_0 <= 27'h0; // @[DCacheMSHR.scala 51:33]
    end else if (!(missReq_fire & secondary_miss)) begin // @[DCacheMSHR.scala 147:39]
      if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
        if (2'h0 == entryStatus_io_next) begin // @[DCacheMSHR.scala 150:43]
          blockAddr_Access_0 <= io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 150:43]
        end
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 51:33]
      blockAddr_Access_1 <= 27'h0; // @[DCacheMSHR.scala 51:33]
    end else if (!(missReq_fire & secondary_miss)) begin // @[DCacheMSHR.scala 147:39]
      if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
        if (2'h1 == entryStatus_io_next) begin // @[DCacheMSHR.scala 150:43]
          blockAddr_Access_1 <= io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 150:43]
        end
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 51:33]
      blockAddr_Access_2 <= 27'h0; // @[DCacheMSHR.scala 51:33]
    end else if (!(missReq_fire & secondary_miss)) begin // @[DCacheMSHR.scala 147:39]
      if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
        if (2'h2 == entryStatus_io_next) begin // @[DCacheMSHR.scala 150:43]
          blockAddr_Access_2 <= io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 150:43]
        end
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 51:33]
      blockAddr_Access_3 <= 27'h0; // @[DCacheMSHR.scala 51:33]
    end else if (!(missReq_fire & secondary_miss)) begin // @[DCacheMSHR.scala 147:39]
      if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
        if (2'h3 == entryStatus_io_next) begin // @[DCacheMSHR.scala 150:43]
          blockAddr_Access_3 <= io_missReq_bits_blockAddr; // @[DCacheMSHR.scala 150:43]
        end
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_0_0 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h0 == _real_SRAMAddrUp_T_3 & _T_58) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_0_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end else if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
      if (2'h0 == entryStatus_io_next) begin // @[DCacheMSHR.scala 151:46]
        instrId_Access_0_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 151:46]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_0_1 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h0 == _real_SRAMAddrUp_T_3 & _T_74) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_0_1 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_0_2 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h0 == _real_SRAMAddrUp_T_3 & _T_90) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_0_2 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_0_3 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h0 == _real_SRAMAddrUp_T_3 & _T_106) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_0_3 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_1_0 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h1 == _real_SRAMAddrUp_T_3 & _T_58) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_1_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end else if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
      if (2'h1 == entryStatus_io_next) begin // @[DCacheMSHR.scala 151:46]
        instrId_Access_1_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 151:46]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_1_1 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h1 == _real_SRAMAddrUp_T_3 & _T_74) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_1_1 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_1_2 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h1 == _real_SRAMAddrUp_T_3 & _T_90) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_1_2 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_1_3 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h1 == _real_SRAMAddrUp_T_3 & _T_106) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_1_3 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_2_0 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h2 == _real_SRAMAddrUp_T_3 & _T_58) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_2_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end else if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
      if (2'h2 == entryStatus_io_next) begin // @[DCacheMSHR.scala 151:46]
        instrId_Access_2_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 151:46]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_2_1 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h2 == _real_SRAMAddrUp_T_3 & _T_74) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_2_1 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_2_2 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h2 == _real_SRAMAddrUp_T_3 & _T_90) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_2_2 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_2_3 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h2 == _real_SRAMAddrUp_T_3 & _T_106) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_2_3 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_3_0 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h3 == _real_SRAMAddrUp_T_3 & _T_58) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_3_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end else if (missReq_fire & primary_miss) begin // @[DCacheMSHR.scala 149:43]
      if (2'h3 == entryStatus_io_next) begin // @[DCacheMSHR.scala 151:46]
        instrId_Access_3_0 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 151:46]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_3_1 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h3 == _real_SRAMAddrUp_T_3 & _T_74) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_3_1 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_3_2 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h3 == _real_SRAMAddrUp_T_3 & _T_90) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_3_2 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 52:31]
      instrId_Access_3_3 <= 2'h0; // @[DCacheMSHR.scala 52:31]
    end else if (missReq_fire & secondary_miss) begin // @[DCacheMSHR.scala 147:39]
      if (2'h3 == _real_SRAMAddrUp_T_3 & _T_106) begin // @[DCacheMSHR.scala 148:73]
        instrId_Access_3_3 <= io_missReq_bits_instrId; // @[DCacheMSHR.scala 148:73]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_0_0 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h0 == real_SRAMAddrUp & 2'h0 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_0_0 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_0_1 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h0 == real_SRAMAddrUp & 2'h1 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_0_1 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_0_2 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h0 == real_SRAMAddrUp & 2'h2 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_0_2 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_0_3 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h0 == real_SRAMAddrUp & 2'h3 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_0_3 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_1_0 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h1 == real_SRAMAddrUp & 2'h0 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_1_0 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_1_1 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h1 == real_SRAMAddrUp & 2'h1 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_1_1 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_1_2 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h1 == real_SRAMAddrUp & 2'h2 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_1_2 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_1_3 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h1 == real_SRAMAddrUp & 2'h3 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_1_3 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_2_0 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h2 == real_SRAMAddrUp & 2'h0 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_2_0 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_2_1 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h2 == real_SRAMAddrUp & 2'h1 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_2_1 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_2_2 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h2 == real_SRAMAddrUp & 2'h2 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_2_2 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_2_3 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h2 == real_SRAMAddrUp & 2'h3 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_2_3 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_3_0 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h3 == real_SRAMAddrUp & 2'h0 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_3_0 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_3_1 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h3 == real_SRAMAddrUp & 2'h1 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_3_1 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_3_2 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h3 == real_SRAMAddrUp & 2'h2 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_3_2 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 53:35]
      targetInfo_Accesss_3_3 <= 65'h0; // @[DCacheMSHR.scala 53:35]
    end else if (missReq_fire) begin // @[DCacheMSHR.scala 105:22]
      if (2'h3 == real_SRAMAddrUp & 2'h3 == real_SRAMAddrDown) begin // @[DCacheMSHR.scala 106:60]
        targetInfo_Accesss_3_3 <= io_missReq_bits_targetInfo; // @[DCacheMSHR.scala 106:60]
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_0_0 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else begin
      subentry_valid_0_0 <= _GEN_73;
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_0_1 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_252) begin // @[DCacheMSHR.scala 135:61]
      if (_T_73) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_0_1 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_0_1 <= _GEN_74;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_0_2 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_252) begin // @[DCacheMSHR.scala 135:61]
      if (_T_89) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_0_2 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_0_2 <= _GEN_78;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_0_3 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_252) begin // @[DCacheMSHR.scala 135:61]
      if (_T_105) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_0_3 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_0_3 <= _GEN_82;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_1_0 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else begin
      subentry_valid_1_0 <= _GEN_89;
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_1_1 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_258) begin // @[DCacheMSHR.scala 135:61]
      if (_T_73) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_1_1 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_1_1 <= _GEN_90;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_1_2 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_258) begin // @[DCacheMSHR.scala 135:61]
      if (_T_89) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_1_2 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_1_2 <= _GEN_94;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_1_3 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_258) begin // @[DCacheMSHR.scala 135:61]
      if (_T_105) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_1_3 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_1_3 <= _GEN_98;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_2_0 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else begin
      subentry_valid_2_0 <= _GEN_105;
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_2_1 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_266) begin // @[DCacheMSHR.scala 135:61]
      if (_T_73) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_2_1 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_2_1 <= _GEN_106;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_2_2 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_266) begin // @[DCacheMSHR.scala 135:61]
      if (_T_89) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_2_2 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_2_2 <= _GEN_110;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_2_3 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_266) begin // @[DCacheMSHR.scala 135:61]
      if (_T_105) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_2_3 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_2_3 <= _GEN_114;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_3_0 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else begin
      subentry_valid_3_0 <= _GEN_121;
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_3_1 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_274) begin // @[DCacheMSHR.scala 135:61]
      if (_T_73) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_3_1 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_3_1 <= _GEN_122;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_3_2 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_274) begin // @[DCacheMSHR.scala 135:61]
      if (_T_89) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_3_2 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_3_2 <= _GEN_126;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 75:31]
      subentry_valid_3_3 <= 1'h0; // @[DCacheMSHR.scala 75:31]
    end else if (_GEN_274) begin // @[DCacheMSHR.scala 135:61]
      if (_T_105) begin // @[DCacheMSHR.scala 137:32]
        subentry_valid_3_3 <= 1'h0; // @[DCacheMSHR.scala 138:43]
      end else begin
        subentry_valid_3_3 <= _GEN_130;
      end
    end
    if (reset) begin // @[DCacheMSHR.scala 96:28]
      missRspBusy <= 1'h0; // @[DCacheMSHR.scala 96:28]
    end else begin
      missRspBusy <= _GEN_49;
    end
    if (reset) begin // @[DCacheMSHR.scala 155:29]
      has_send2mem_0 <= 1'h0; // @[DCacheMSHR.scala 155:29]
    end else begin
      has_send2mem_0 <= _GEN_199;
    end
    if (reset) begin // @[DCacheMSHR.scala 155:29]
      has_send2mem_1 <= 1'h0; // @[DCacheMSHR.scala 155:29]
    end else begin
      has_send2mem_1 <= _GEN_193;
    end
    if (reset) begin // @[DCacheMSHR.scala 155:29]
      has_send2mem_2 <= 1'h0; // @[DCacheMSHR.scala 155:29]
    end else begin
      has_send2mem_2 <= _GEN_195;
    end
    if (reset) begin // @[DCacheMSHR.scala 155:29]
      has_send2mem_3 <= 1'h0; // @[DCacheMSHR.scala 155:29]
    end else begin
      has_send2mem_3 <= _GEN_197;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(_T_8 <= 3'h1)) begin
          $fatal; // @[DCacheMSHR.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_8 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCacheMSHR.scala:88 assert(PopCount(entryMatchMissRsp) <= 1.U)\n"); // @[DCacheMSHR.scala 88:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_12 & ~(_T_22 <= 3'h1)) begin
          $fatal; // @[DCacheMSHR.scala 90:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_12 & ~(_T_22 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCacheMSHR.scala:90 assert(PopCount(entryMatchMissReq) <= 1.U)\n"); // @[DCacheMSHR.scala 90:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_12 & ~(~_T_28 | _T_28 & subentryStatus_io_used >= 3'h1)) begin
          $fatal; // @[DCacheMSHR.scala 115:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_12 & ~(~_T_28 | _T_28 & subentryStatus_io_used >= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCacheMSHR.scala:115 assert(!io.missRspIn.fire || (io.missRspIn.fire && subentryStatus.io.used >= 1.U))\n"
            ); // @[DCacheMSHR.scala 115:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  blockAddr_Access_0 = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  blockAddr_Access_1 = _RAND_1[26:0];
  _RAND_2 = {1{`RANDOM}};
  blockAddr_Access_2 = _RAND_2[26:0];
  _RAND_3 = {1{`RANDOM}};
  blockAddr_Access_3 = _RAND_3[26:0];
  _RAND_4 = {1{`RANDOM}};
  instrId_Access_0_0 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  instrId_Access_0_1 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  instrId_Access_0_2 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  instrId_Access_0_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  instrId_Access_1_0 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  instrId_Access_1_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  instrId_Access_1_2 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  instrId_Access_1_3 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  instrId_Access_2_0 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  instrId_Access_2_1 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  instrId_Access_2_2 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  instrId_Access_2_3 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  instrId_Access_3_0 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  instrId_Access_3_1 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  instrId_Access_3_2 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  instrId_Access_3_3 = _RAND_19[1:0];
  _RAND_20 = {3{`RANDOM}};
  targetInfo_Accesss_0_0 = _RAND_20[64:0];
  _RAND_21 = {3{`RANDOM}};
  targetInfo_Accesss_0_1 = _RAND_21[64:0];
  _RAND_22 = {3{`RANDOM}};
  targetInfo_Accesss_0_2 = _RAND_22[64:0];
  _RAND_23 = {3{`RANDOM}};
  targetInfo_Accesss_0_3 = _RAND_23[64:0];
  _RAND_24 = {3{`RANDOM}};
  targetInfo_Accesss_1_0 = _RAND_24[64:0];
  _RAND_25 = {3{`RANDOM}};
  targetInfo_Accesss_1_1 = _RAND_25[64:0];
  _RAND_26 = {3{`RANDOM}};
  targetInfo_Accesss_1_2 = _RAND_26[64:0];
  _RAND_27 = {3{`RANDOM}};
  targetInfo_Accesss_1_3 = _RAND_27[64:0];
  _RAND_28 = {3{`RANDOM}};
  targetInfo_Accesss_2_0 = _RAND_28[64:0];
  _RAND_29 = {3{`RANDOM}};
  targetInfo_Accesss_2_1 = _RAND_29[64:0];
  _RAND_30 = {3{`RANDOM}};
  targetInfo_Accesss_2_2 = _RAND_30[64:0];
  _RAND_31 = {3{`RANDOM}};
  targetInfo_Accesss_2_3 = _RAND_31[64:0];
  _RAND_32 = {3{`RANDOM}};
  targetInfo_Accesss_3_0 = _RAND_32[64:0];
  _RAND_33 = {3{`RANDOM}};
  targetInfo_Accesss_3_1 = _RAND_33[64:0];
  _RAND_34 = {3{`RANDOM}};
  targetInfo_Accesss_3_2 = _RAND_34[64:0];
  _RAND_35 = {3{`RANDOM}};
  targetInfo_Accesss_3_3 = _RAND_35[64:0];
  _RAND_36 = {1{`RANDOM}};
  subentry_valid_0_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  subentry_valid_0_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  subentry_valid_0_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  subentry_valid_0_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  subentry_valid_1_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  subentry_valid_1_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  subentry_valid_1_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  subentry_valid_1_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  subentry_valid_2_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  subentry_valid_2_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  subentry_valid_2_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  subentry_valid_2_3 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  subentry_valid_3_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  subentry_valid_3_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  subentry_valid_3_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  subentry_valid_3_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  missRspBusy = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  has_send2mem_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  has_send2mem_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  has_send2mem_2 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  has_send2mem_3 = _RAND_56[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataCrossbar(
  input  [31:0] io_DataIn_0,
  input  [31:0] io_DataIn_1,
  input  [31:0] io_DataIn_2,
  input  [31:0] io_DataIn_3,
  input  [31:0] io_DataIn_4,
  input  [31:0] io_DataIn_5,
  input  [31:0] io_DataIn_6,
  input  [31:0] io_DataIn_7,
  output [31:0] io_DataOut_0,
  output [31:0] io_DataOut_1,
  output [31:0] io_DataOut_2,
  output [31:0] io_DataOut_3,
  output [31:0] io_DataOut_4,
  output [31:0] io_DataOut_5,
  output [31:0] io_DataOut_6,
  output [31:0] io_DataOut_7,
  input  [7:0]  io_Select1H_0,
  input  [7:0]  io_Select1H_1,
  input  [7:0]  io_Select1H_2,
  input  [7:0]  io_Select1H_3,
  input  [7:0]  io_Select1H_4,
  input  [7:0]  io_Select1H_5,
  input  [7:0]  io_Select1H_6,
  input  [7:0]  io_Select1H_7
);
  wire [31:0] _io_DataOut_0_T_8 = io_Select1H_0[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_9 = io_Select1H_0[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_10 = io_Select1H_0[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_11 = io_Select1H_0[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_12 = io_Select1H_0[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_13 = io_Select1H_0[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_14 = io_Select1H_0[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_15 = io_Select1H_0[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_16 = _io_DataOut_0_T_8 | _io_DataOut_0_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_17 = _io_DataOut_0_T_16 | _io_DataOut_0_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_18 = _io_DataOut_0_T_17 | _io_DataOut_0_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_19 = _io_DataOut_0_T_18 | _io_DataOut_0_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_20 = _io_DataOut_0_T_19 | _io_DataOut_0_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_0_T_21 = _io_DataOut_0_T_20 | _io_DataOut_0_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_8 = io_Select1H_1[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_9 = io_Select1H_1[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_10 = io_Select1H_1[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_11 = io_Select1H_1[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_12 = io_Select1H_1[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_13 = io_Select1H_1[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_14 = io_Select1H_1[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_15 = io_Select1H_1[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_16 = _io_DataOut_1_T_8 | _io_DataOut_1_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_17 = _io_DataOut_1_T_16 | _io_DataOut_1_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_18 = _io_DataOut_1_T_17 | _io_DataOut_1_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_19 = _io_DataOut_1_T_18 | _io_DataOut_1_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_20 = _io_DataOut_1_T_19 | _io_DataOut_1_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_1_T_21 = _io_DataOut_1_T_20 | _io_DataOut_1_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_8 = io_Select1H_2[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_9 = io_Select1H_2[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_10 = io_Select1H_2[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_11 = io_Select1H_2[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_12 = io_Select1H_2[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_13 = io_Select1H_2[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_14 = io_Select1H_2[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_15 = io_Select1H_2[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_16 = _io_DataOut_2_T_8 | _io_DataOut_2_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_17 = _io_DataOut_2_T_16 | _io_DataOut_2_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_18 = _io_DataOut_2_T_17 | _io_DataOut_2_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_19 = _io_DataOut_2_T_18 | _io_DataOut_2_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_20 = _io_DataOut_2_T_19 | _io_DataOut_2_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_2_T_21 = _io_DataOut_2_T_20 | _io_DataOut_2_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_8 = io_Select1H_3[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_9 = io_Select1H_3[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_10 = io_Select1H_3[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_11 = io_Select1H_3[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_12 = io_Select1H_3[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_13 = io_Select1H_3[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_14 = io_Select1H_3[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_15 = io_Select1H_3[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_16 = _io_DataOut_3_T_8 | _io_DataOut_3_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_17 = _io_DataOut_3_T_16 | _io_DataOut_3_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_18 = _io_DataOut_3_T_17 | _io_DataOut_3_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_19 = _io_DataOut_3_T_18 | _io_DataOut_3_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_20 = _io_DataOut_3_T_19 | _io_DataOut_3_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_3_T_21 = _io_DataOut_3_T_20 | _io_DataOut_3_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_8 = io_Select1H_4[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_9 = io_Select1H_4[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_10 = io_Select1H_4[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_11 = io_Select1H_4[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_12 = io_Select1H_4[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_13 = io_Select1H_4[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_14 = io_Select1H_4[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_15 = io_Select1H_4[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_16 = _io_DataOut_4_T_8 | _io_DataOut_4_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_17 = _io_DataOut_4_T_16 | _io_DataOut_4_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_18 = _io_DataOut_4_T_17 | _io_DataOut_4_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_19 = _io_DataOut_4_T_18 | _io_DataOut_4_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_20 = _io_DataOut_4_T_19 | _io_DataOut_4_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_4_T_21 = _io_DataOut_4_T_20 | _io_DataOut_4_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_8 = io_Select1H_5[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_9 = io_Select1H_5[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_10 = io_Select1H_5[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_11 = io_Select1H_5[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_12 = io_Select1H_5[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_13 = io_Select1H_5[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_14 = io_Select1H_5[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_15 = io_Select1H_5[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_16 = _io_DataOut_5_T_8 | _io_DataOut_5_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_17 = _io_DataOut_5_T_16 | _io_DataOut_5_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_18 = _io_DataOut_5_T_17 | _io_DataOut_5_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_19 = _io_DataOut_5_T_18 | _io_DataOut_5_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_20 = _io_DataOut_5_T_19 | _io_DataOut_5_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_5_T_21 = _io_DataOut_5_T_20 | _io_DataOut_5_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_8 = io_Select1H_6[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_9 = io_Select1H_6[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_10 = io_Select1H_6[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_11 = io_Select1H_6[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_12 = io_Select1H_6[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_13 = io_Select1H_6[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_14 = io_Select1H_6[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_15 = io_Select1H_6[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_16 = _io_DataOut_6_T_8 | _io_DataOut_6_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_17 = _io_DataOut_6_T_16 | _io_DataOut_6_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_18 = _io_DataOut_6_T_17 | _io_DataOut_6_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_19 = _io_DataOut_6_T_18 | _io_DataOut_6_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_20 = _io_DataOut_6_T_19 | _io_DataOut_6_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_6_T_21 = _io_DataOut_6_T_20 | _io_DataOut_6_T_14; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_8 = io_Select1H_7[0] ? io_DataIn_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_9 = io_Select1H_7[1] ? io_DataIn_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_10 = io_Select1H_7[2] ? io_DataIn_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_11 = io_Select1H_7[3] ? io_DataIn_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_12 = io_Select1H_7[4] ? io_DataIn_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_13 = io_Select1H_7[5] ? io_DataIn_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_14 = io_Select1H_7[6] ? io_DataIn_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_15 = io_Select1H_7[7] ? io_DataIn_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_16 = _io_DataOut_7_T_8 | _io_DataOut_7_T_9; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_17 = _io_DataOut_7_T_16 | _io_DataOut_7_T_10; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_18 = _io_DataOut_7_T_17 | _io_DataOut_7_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_19 = _io_DataOut_7_T_18 | _io_DataOut_7_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_20 = _io_DataOut_7_T_19 | _io_DataOut_7_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_DataOut_7_T_21 = _io_DataOut_7_T_20 | _io_DataOut_7_T_14; // @[Mux.scala 27:73]
  assign io_DataOut_0 = _io_DataOut_0_T_21 | _io_DataOut_0_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_1 = _io_DataOut_1_T_21 | _io_DataOut_1_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_2 = _io_DataOut_2_T_21 | _io_DataOut_2_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_3 = _io_DataOut_3_T_21 | _io_DataOut_3_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_4 = _io_DataOut_4_T_21 | _io_DataOut_4_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_5 = _io_DataOut_5_T_21 | _io_DataOut_5_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_6 = _io_DataOut_6_T_21 | _io_DataOut_6_T_15; // @[Mux.scala 27:73]
  assign io_DataOut_7 = _io_DataOut_7_T_21 | _io_DataOut_7_T_15; // @[Mux.scala 27:73]
endmodule
module WdbEnqPtrGen(
  input        io_entryValidList_0,
  input        io_entryValidList_1,
  input        io_entryValidList_2,
  input        io_entryValidList_3,
  input  [1:0] io_enqPtr_cs,
  output [1:0] io_enqPtr_ns
);
  wire [2:0] _muxSel_T = {{1'd0}, io_enqPtr_cs}; // @[WDB.scala 42:19]
  wire [1:0] muxSel = _muxSel_T[1:0] + 2'h1; // @[WDB.scala 42:34]
  wire [3:0] _cyclicValidList_0_T = 4'h1 << muxSel; // @[OneHot.scala 57:35]
  wire  cyclicValidList_0 = _cyclicValidList_0_T[0] & io_entryValidList_0 | _cyclicValidList_0_T[1] &
    io_entryValidList_1 | _cyclicValidList_0_T[2] & io_entryValidList_2 | _cyclicValidList_0_T[3] & io_entryValidList_3; // @[Mux.scala 27:73]
  wire [1:0] _muxSel_T_5 = 2'h1 + io_enqPtr_cs; // @[WDB.scala 42:19]
  wire [1:0] muxSel_1 = _muxSel_T_5 + 2'h1; // @[WDB.scala 42:34]
  wire [3:0] _cyclicValidList_1_T = 4'h1 << muxSel_1; // @[OneHot.scala 57:35]
  wire  cyclicValidList_1 = _cyclicValidList_1_T[0] & io_entryValidList_0 | _cyclicValidList_1_T[1] &
    io_entryValidList_1 | _cyclicValidList_1_T[2] & io_entryValidList_2 | _cyclicValidList_1_T[3] & io_entryValidList_3; // @[Mux.scala 27:73]
  wire [1:0] _muxSel_T_9 = 2'h2 + io_enqPtr_cs; // @[WDB.scala 42:19]
  wire [1:0] muxSel_2 = _muxSel_T_9 + 2'h1; // @[WDB.scala 42:34]
  wire [3:0] _cyclicValidList_2_T = 4'h1 << muxSel_2; // @[OneHot.scala 57:35]
  wire  cyclicValidList_2 = _cyclicValidList_2_T[0] & io_entryValidList_0 | _cyclicValidList_2_T[1] &
    io_entryValidList_1 | _cyclicValidList_2_T[2] & io_entryValidList_2 | _cyclicValidList_2_T[3] & io_entryValidList_3; // @[Mux.scala 27:73]
  wire  _io_enqPtr_ns_T = ~cyclicValidList_0; // @[WDB.scala 45:55]
  wire  _io_enqPtr_ns_T_1 = ~cyclicValidList_1; // @[WDB.scala 45:55]
  wire  _io_enqPtr_ns_T_2 = ~cyclicValidList_2; // @[WDB.scala 45:55]
  wire [1:0] _io_enqPtr_ns_T_4 = _io_enqPtr_ns_T_2 ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _io_enqPtr_ns_T_5 = _io_enqPtr_ns_T_1 ? 2'h1 : _io_enqPtr_ns_T_4; // @[Mux.scala 47:70]
  wire [1:0] _io_enqPtr_ns_T_6 = _io_enqPtr_ns_T ? 2'h0 : _io_enqPtr_ns_T_5; // @[Mux.scala 47:70]
  wire [1:0] _io_enqPtr_ns_T_8 = _io_enqPtr_ns_T_6 + 2'h1; // @[WDB.scala 45:60]
  assign io_enqPtr_ns = _io_enqPtr_ns_T_8 + io_enqPtr_cs; // @[WDB.scala 45:66]
endmodule
module WdbDeqPtrGen(
  input        io_entryValidList_0,
  input        io_entryValidList_1,
  input        io_entryValidList_2,
  input        io_entryValidList_3,
  input        io_entryFrozenList_0,
  input        io_entryFrozenList_1,
  input        io_entryFrozenList_2,
  input        io_entryFrozenList_3,
  input  [1:0] io_deqPtr_cs,
  output [1:0] io_deqPtr_ns
);
  wire [3:0] _UnfrozenValidList_T = {io_entryValidList_0,io_entryValidList_1,io_entryValidList_2,io_entryValidList_3}; // @[Cat.scala 31:58]
  wire [3:0] _UnfrozenValidList_T_1 = {io_entryFrozenList_0,io_entryFrozenList_1,io_entryFrozenList_2,
    io_entryFrozenList_3}; // @[Cat.scala 31:58]
  wire [3:0] _UnfrozenValidList_T_2 = _UnfrozenValidList_T ^ _UnfrozenValidList_T_1; // @[WDB.scala 71:58]
  wire [3:0] UnfrozenValidList = {_UnfrozenValidList_T_2[0],_UnfrozenValidList_T_2[1],_UnfrozenValidList_T_2[2],
    _UnfrozenValidList_T_2[3]}; // @[Cat.scala 31:58]
  wire [2:0] _muxSel_T = {{1'd0}, io_deqPtr_cs}; // @[WDB.scala 76:19]
  wire [1:0] muxSel = _muxSel_T[1:0] + 2'h1; // @[WDB.scala 76:34]
  wire [3:0] _cyclicValidList_0_T = 4'h1 << muxSel; // @[OneHot.scala 57:35]
  wire [3:0] _cyclicValidList_0_T_1 = _cyclicValidList_0_T & UnfrozenValidList; // @[Mux.scala 30:47]
  wire  cyclicValidList_0 = |_cyclicValidList_0_T_1; // @[Mux.scala 30:53]
  wire [1:0] _muxSel_T_5 = 2'h1 + io_deqPtr_cs; // @[WDB.scala 76:19]
  wire [1:0] muxSel_1 = _muxSel_T_5 + 2'h1; // @[WDB.scala 76:34]
  wire [3:0] _cyclicValidList_1_T = 4'h1 << muxSel_1; // @[OneHot.scala 57:35]
  wire [3:0] _cyclicValidList_1_T_1 = _cyclicValidList_1_T & UnfrozenValidList; // @[Mux.scala 30:47]
  wire  cyclicValidList_1 = |_cyclicValidList_1_T_1; // @[Mux.scala 30:53]
  wire [1:0] _muxSel_T_9 = 2'h2 + io_deqPtr_cs; // @[WDB.scala 76:19]
  wire [1:0] muxSel_2 = _muxSel_T_9 + 2'h1; // @[WDB.scala 76:34]
  wire [3:0] _cyclicValidList_2_T = 4'h1 << muxSel_2; // @[OneHot.scala 57:35]
  wire [3:0] _cyclicValidList_2_T_1 = _cyclicValidList_2_T & UnfrozenValidList; // @[Mux.scala 30:47]
  wire  cyclicValidList_2 = |_cyclicValidList_2_T_1; // @[Mux.scala 30:53]
  wire [1:0] _io_deqPtr_ns_T = cyclicValidList_2 ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _io_deqPtr_ns_T_1 = cyclicValidList_1 ? 2'h1 : _io_deqPtr_ns_T; // @[Mux.scala 47:70]
  wire [1:0] _io_deqPtr_ns_T_2 = cyclicValidList_0 ? 2'h0 : _io_deqPtr_ns_T_1; // @[Mux.scala 47:70]
  wire [1:0] _io_deqPtr_ns_T_4 = _io_deqPtr_ns_T_2 + 2'h1; // @[WDB.scala 80:52]
  assign io_deqPtr_ns = _io_deqPtr_ns_T_4 + io_deqPtr_cs; // @[WDB.scala 80:58]
endmodule
module WDB(
  input         clock,
  input         reset,
  output        io_inputBus_ready,
  input         io_inputBus_valid,
  input  [3:0]  io_inputBus_bits_mask_0,
  input  [3:0]  io_inputBus_bits_mask_1,
  input  [3:0]  io_inputBus_bits_mask_2,
  input  [3:0]  io_inputBus_bits_mask_3,
  input  [3:0]  io_inputBus_bits_mask_4,
  input  [3:0]  io_inputBus_bits_mask_5,
  input  [3:0]  io_inputBus_bits_mask_6,
  input  [3:0]  io_inputBus_bits_mask_7,
  input  [31:0] io_inputBus_bits_addr,
  input  [7:0]  io_inputBus_bits_data_0_0,
  input  [7:0]  io_inputBus_bits_data_0_1,
  input  [7:0]  io_inputBus_bits_data_0_2,
  input  [7:0]  io_inputBus_bits_data_0_3,
  input  [7:0]  io_inputBus_bits_data_1_0,
  input  [7:0]  io_inputBus_bits_data_1_1,
  input  [7:0]  io_inputBus_bits_data_1_2,
  input  [7:0]  io_inputBus_bits_data_1_3,
  input  [7:0]  io_inputBus_bits_data_2_0,
  input  [7:0]  io_inputBus_bits_data_2_1,
  input  [7:0]  io_inputBus_bits_data_2_2,
  input  [7:0]  io_inputBus_bits_data_2_3,
  input  [7:0]  io_inputBus_bits_data_3_0,
  input  [7:0]  io_inputBus_bits_data_3_1,
  input  [7:0]  io_inputBus_bits_data_3_2,
  input  [7:0]  io_inputBus_bits_data_3_3,
  input  [7:0]  io_inputBus_bits_data_4_0,
  input  [7:0]  io_inputBus_bits_data_4_1,
  input  [7:0]  io_inputBus_bits_data_4_2,
  input  [7:0]  io_inputBus_bits_data_4_3,
  input  [7:0]  io_inputBus_bits_data_5_0,
  input  [7:0]  io_inputBus_bits_data_5_1,
  input  [7:0]  io_inputBus_bits_data_5_2,
  input  [7:0]  io_inputBus_bits_data_5_3,
  input  [7:0]  io_inputBus_bits_data_6_0,
  input  [7:0]  io_inputBus_bits_data_6_1,
  input  [7:0]  io_inputBus_bits_data_6_2,
  input  [7:0]  io_inputBus_bits_data_6_3,
  input  [7:0]  io_inputBus_bits_data_7_0,
  input  [7:0]  io_inputBus_bits_data_7_1,
  input  [7:0]  io_inputBus_bits_data_7_2,
  input  [7:0]  io_inputBus_bits_data_7_3,
  input  [1:0]  io_inputBus_bits_instrId,
  input         io_inputBus_bits_bankConflict,
  input         io_inputBus_bits_subWordMissReq,
  input         io_inputBus_bits_subWordMissRsp,
  input         io_outputBus_ready,
  output        io_outputBus_valid,
  output        io_outputBus_bits_mask_0,
  output        io_outputBus_bits_mask_1,
  output        io_outputBus_bits_mask_2,
  output        io_outputBus_bits_mask_3,
  output        io_outputBus_bits_mask_4,
  output        io_outputBus_bits_mask_5,
  output        io_outputBus_bits_mask_6,
  output        io_outputBus_bits_mask_7,
  output [31:0] io_outputBus_bits_addr,
  output [7:0]  io_outputBus_bits_data_0_0,
  output [7:0]  io_outputBus_bits_data_0_1,
  output [7:0]  io_outputBus_bits_data_0_2,
  output [7:0]  io_outputBus_bits_data_0_3,
  output [7:0]  io_outputBus_bits_data_1_0,
  output [7:0]  io_outputBus_bits_data_1_1,
  output [7:0]  io_outputBus_bits_data_1_2,
  output [7:0]  io_outputBus_bits_data_1_3,
  output [7:0]  io_outputBus_bits_data_2_0,
  output [7:0]  io_outputBus_bits_data_2_1,
  output [7:0]  io_outputBus_bits_data_2_2,
  output [7:0]  io_outputBus_bits_data_2_3,
  output [7:0]  io_outputBus_bits_data_3_0,
  output [7:0]  io_outputBus_bits_data_3_1,
  output [7:0]  io_outputBus_bits_data_3_2,
  output [7:0]  io_outputBus_bits_data_3_3,
  output [7:0]  io_outputBus_bits_data_4_0,
  output [7:0]  io_outputBus_bits_data_4_1,
  output [7:0]  io_outputBus_bits_data_4_2,
  output [7:0]  io_outputBus_bits_data_4_3,
  output [7:0]  io_outputBus_bits_data_5_0,
  output [7:0]  io_outputBus_bits_data_5_1,
  output [7:0]  io_outputBus_bits_data_5_2,
  output [7:0]  io_outputBus_bits_data_5_3,
  output [7:0]  io_outputBus_bits_data_6_0,
  output [7:0]  io_outputBus_bits_data_6_1,
  output [7:0]  io_outputBus_bits_data_6_2,
  output [7:0]  io_outputBus_bits_data_6_3,
  output [7:0]  io_outputBus_bits_data_7_0,
  output [7:0]  io_outputBus_bits_data_7_1,
  output [7:0]  io_outputBus_bits_data_7_2,
  output [7:0]  io_outputBus_bits_data_7_3,
  output [1:0]  io_outputBus_bits_instrId,
  output        io_wdbAlmostFull
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
`endif // RANDOMIZE_REG_INIT
  wire  enqPtr_w_Gen_io_entryValidList_0; // @[WDB.scala 53:21]
  wire  enqPtr_w_Gen_io_entryValidList_1; // @[WDB.scala 53:21]
  wire  enqPtr_w_Gen_io_entryValidList_2; // @[WDB.scala 53:21]
  wire  enqPtr_w_Gen_io_entryValidList_3; // @[WDB.scala 53:21]
  wire [1:0] enqPtr_w_Gen_io_enqPtr_cs; // @[WDB.scala 53:21]
  wire [1:0] enqPtr_w_Gen_io_enqPtr_ns; // @[WDB.scala 53:21]
  wire  deqPtr_w_Gen_io_entryValidList_0; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryValidList_1; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryValidList_2; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryValidList_3; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryFrozenList_0; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryFrozenList_1; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryFrozenList_2; // @[WDB.scala 89:21]
  wire  deqPtr_w_Gen_io_entryFrozenList_3; // @[WDB.scala 89:21]
  wire [1:0] deqPtr_w_Gen_io_deqPtr_cs; // @[WDB.scala 89:21]
  wire [1:0] deqPtr_w_Gen_io_deqPtr_ns; // @[WDB.scala 89:21]
  reg  mask_ram_0_0; // @[WDB.scala 104:25]
  reg  mask_ram_0_1; // @[WDB.scala 104:25]
  reg  mask_ram_0_2; // @[WDB.scala 104:25]
  reg  mask_ram_0_3; // @[WDB.scala 104:25]
  reg  mask_ram_0_4; // @[WDB.scala 104:25]
  reg  mask_ram_0_5; // @[WDB.scala 104:25]
  reg  mask_ram_0_6; // @[WDB.scala 104:25]
  reg  mask_ram_0_7; // @[WDB.scala 104:25]
  reg  mask_ram_1_0; // @[WDB.scala 104:25]
  reg  mask_ram_1_1; // @[WDB.scala 104:25]
  reg  mask_ram_1_2; // @[WDB.scala 104:25]
  reg  mask_ram_1_3; // @[WDB.scala 104:25]
  reg  mask_ram_1_4; // @[WDB.scala 104:25]
  reg  mask_ram_1_5; // @[WDB.scala 104:25]
  reg  mask_ram_1_6; // @[WDB.scala 104:25]
  reg  mask_ram_1_7; // @[WDB.scala 104:25]
  reg  mask_ram_2_0; // @[WDB.scala 104:25]
  reg  mask_ram_2_1; // @[WDB.scala 104:25]
  reg  mask_ram_2_2; // @[WDB.scala 104:25]
  reg  mask_ram_2_3; // @[WDB.scala 104:25]
  reg  mask_ram_2_4; // @[WDB.scala 104:25]
  reg  mask_ram_2_5; // @[WDB.scala 104:25]
  reg  mask_ram_2_6; // @[WDB.scala 104:25]
  reg  mask_ram_2_7; // @[WDB.scala 104:25]
  reg  mask_ram_3_0; // @[WDB.scala 104:25]
  reg  mask_ram_3_1; // @[WDB.scala 104:25]
  reg  mask_ram_3_2; // @[WDB.scala 104:25]
  reg  mask_ram_3_3; // @[WDB.scala 104:25]
  reg  mask_ram_3_4; // @[WDB.scala 104:25]
  reg  mask_ram_3_5; // @[WDB.scala 104:25]
  reg  mask_ram_3_6; // @[WDB.scala 104:25]
  reg  mask_ram_3_7; // @[WDB.scala 104:25]
  reg [31:0] addr_ram_0; // @[WDB.scala 105:25]
  reg [31:0] addr_ram_1; // @[WDB.scala 105:25]
  reg [31:0] addr_ram_2; // @[WDB.scala 105:25]
  reg [31:0] addr_ram_3; // @[WDB.scala 105:25]
  reg [7:0] data_ram_0_0_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_0_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_0_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_0_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_1_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_1_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_1_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_1_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_2_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_2_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_2_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_2_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_3_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_3_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_3_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_3_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_4_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_4_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_4_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_4_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_5_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_5_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_5_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_5_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_6_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_6_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_6_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_6_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_7_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_7_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_7_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_0_7_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_0_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_0_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_0_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_0_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_1_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_1_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_1_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_1_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_2_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_2_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_2_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_2_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_3_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_3_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_3_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_3_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_4_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_4_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_4_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_4_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_5_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_5_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_5_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_5_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_6_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_6_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_6_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_6_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_7_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_7_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_7_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_1_7_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_0_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_0_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_0_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_0_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_1_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_1_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_1_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_1_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_2_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_2_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_2_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_2_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_3_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_3_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_3_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_3_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_4_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_4_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_4_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_4_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_5_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_5_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_5_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_5_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_6_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_6_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_6_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_6_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_7_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_7_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_7_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_2_7_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_0_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_0_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_0_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_0_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_1_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_1_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_1_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_1_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_2_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_2_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_2_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_2_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_3_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_3_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_3_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_3_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_4_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_4_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_4_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_4_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_5_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_5_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_5_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_5_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_6_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_6_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_6_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_6_3; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_7_0; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_7_1; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_7_2; // @[WDB.scala 106:25]
  reg [7:0] data_ram_3_7_3; // @[WDB.scala 106:25]
  reg [1:0] instrId_ram_0; // @[WDB.scala 109:28]
  reg [1:0] instrId_ram_1; // @[WDB.scala 109:28]
  reg [1:0] instrId_ram_2; // @[WDB.scala 109:28]
  reg [1:0] instrId_ram_3; // @[WDB.scala 109:28]
  reg [1:0] enqPtr; // @[WDB.scala 111:23]
  reg [1:0] deqPtr; // @[WDB.scala 112:23]
  reg  entryValid_0; // @[WDB.scala 118:27]
  reg  entryValid_1; // @[WDB.scala 118:27]
  reg  entryValid_2; // @[WDB.scala 118:27]
  reg  entryValid_3; // @[WDB.scala 118:27]
  reg  entryFrozen_0; // @[WDB.scala 119:28]
  reg  entryFrozen_1; // @[WDB.scala 119:28]
  reg  entryFrozen_2; // @[WDB.scala 119:28]
  reg  entryFrozen_3; // @[WDB.scala 119:28]
  wire  doEnq = io_inputBus_ready & io_inputBus_valid; // @[Decoupled.scala 50:35]
  wire  doDeq = io_outputBus_ready & io_outputBus_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _almFull_T = {entryValid_0,entryValid_1,entryValid_2,entryValid_3}; // @[Cat.scala 31:58]
  wire [1:0] _almFull_T_5 = _almFull_T[0] + _almFull_T[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _almFull_T_7 = _almFull_T[2] + _almFull_T[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _almFull_T_9 = _almFull_T_5 + _almFull_T_7; // @[Bitwise.scala 48:55]
  wire  _T_1 = doEnq & ~io_inputBus_bits_bankConflict; // @[WDB.scala 133:15]
  wire [1:0] enqPtr_w = enqPtr_w_Gen_io_enqPtr_ns; // @[WDB.scala 114:22 132:12]
  wire [1:0] deqPtr_w = deqPtr_w_Gen_io_deqPtr_ns; // @[WDB.scala 115:22 137:12]
  wire  meltMatch_0 = addr_ram_0 == io_inputBus_bits_addr; // @[WDB.scala 144:33]
  wire  meltMatch_1 = addr_ram_1 == io_inputBus_bits_addr; // @[WDB.scala 144:33]
  wire  meltMatch_2 = addr_ram_2 == io_inputBus_bits_addr; // @[WDB.scala 144:33]
  wire  meltMatch_3 = addr_ram_3 == io_inputBus_bits_addr; // @[WDB.scala 144:33]
  wire [3:0] _T_2 = {meltMatch_0,meltMatch_1,meltMatch_2,meltMatch_3}; // @[Cat.scala 31:58]
  wire [1:0] _T_7 = _T_2[0] + _T_2[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _T_9 = _T_2[2] + _T_2[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _T_11 = _T_7 + _T_9; // @[Bitwise.scala 48:55]
  wire  _T_15 = ~io_inputBus_bits_subWordMissRsp; // @[WDB.scala 146:64]
  wire  _T_18 = ~reset; // @[WDB.scala 146:9]
  wire [3:0] _meltPtr_w_T = {meltMatch_3,meltMatch_2,meltMatch_1,meltMatch_0}; // @[OneHot.scala 22:45]
  wire [1:0] meltPtr_w_hi_1 = _meltPtr_w_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] meltPtr_w_lo_1 = _meltPtr_w_T[1:0]; // @[OneHot.scala 31:18]
  wire  _meltPtr_w_T_1 = |meltPtr_w_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _meltPtr_w_T_2 = meltPtr_w_hi_1 | meltPtr_w_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] meltPtr_w = {_meltPtr_w_T_1,_meltPtr_w_T_2[1]}; // @[Cat.scala 31:58]
  wire  _GEN_3 = 2'h1 == meltPtr_w ? entryFrozen_1 : entryFrozen_0; // @[WDB.scala 148:{33,33}]
  wire  _GEN_4 = 2'h2 == meltPtr_w ? entryFrozen_2 : _GEN_3; // @[WDB.scala 148:{33,33}]
  wire  _GEN_5 = 2'h3 == meltPtr_w ? entryFrozen_3 : _GEN_4; // @[WDB.scala 148:{33,33}]
  wire  _GEN_6 = io_inputBus_bits_subWordMissReq | entryFrozen_0; // @[WDB.scala 119:28 158:32 159:28]
  wire  _GEN_7 = 2'h0 == enqPtr_w | entryValid_0; // @[WDB.scala 118:27 156:37 157:27]
  wire  _GEN_8 = 2'h0 == enqPtr_w ? _GEN_6 : entryFrozen_0; // @[WDB.scala 119:28 156:37]
  wire  _GEN_14 = io_inputBus_bits_subWordMissReq | entryFrozen_1; // @[WDB.scala 119:28 158:32 159:28]
  wire  _GEN_15 = 2'h1 == enqPtr_w | entryValid_1; // @[WDB.scala 118:27 156:37 157:27]
  wire  _GEN_16 = 2'h1 == enqPtr_w ? _GEN_14 : entryFrozen_1; // @[WDB.scala 119:28 156:37]
  wire  _GEN_22 = io_inputBus_bits_subWordMissReq | entryFrozen_2; // @[WDB.scala 119:28 158:32 159:28]
  wire  _GEN_23 = 2'h2 == enqPtr_w | entryValid_2; // @[WDB.scala 118:27 156:37 157:27]
  wire  _GEN_24 = 2'h2 == enqPtr_w ? _GEN_22 : entryFrozen_2; // @[WDB.scala 119:28 156:37]
  wire  _GEN_30 = io_inputBus_bits_subWordMissReq | entryFrozen_3; // @[WDB.scala 119:28 158:32 159:28]
  wire  _GEN_31 = 2'h3 == enqPtr_w | entryValid_3; // @[WDB.scala 118:27 156:37 157:27]
  wire  _GEN_32 = 2'h3 == enqPtr_w ? _GEN_30 : entryFrozen_3; // @[WDB.scala 119:28 156:37]
  wire  _mask_ram_0_T = &io_inputBus_bits_mask_0; // @[WDB.scala 172:69]
  wire  _GEN_38 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_0 : mask_ram_0_0; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_39 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_0 : mask_ram_1_0; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_40 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_0 : mask_ram_2_0; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_41 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_0 : mask_ram_3_0; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_42 = 2'h0 == meltPtr_w ? _mask_ram_0_T : mask_ram_0_0; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_43 = 2'h1 == meltPtr_w ? _mask_ram_0_T : mask_ram_1_0; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_44 = 2'h2 == meltPtr_w ? _mask_ram_0_T : mask_ram_2_0; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_45 = 2'h3 == meltPtr_w ? _mask_ram_0_T : mask_ram_3_0; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_1_T = &io_inputBus_bits_mask_1; // @[WDB.scala 172:69]
  wire  _GEN_58 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_1 : mask_ram_0_1; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_59 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_1 : mask_ram_1_1; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_60 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_1 : mask_ram_2_1; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_61 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_1 : mask_ram_3_1; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_62 = 2'h0 == meltPtr_w ? _mask_ram_1_T : mask_ram_0_1; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_63 = 2'h1 == meltPtr_w ? _mask_ram_1_T : mask_ram_1_1; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_64 = 2'h2 == meltPtr_w ? _mask_ram_1_T : mask_ram_2_1; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_65 = 2'h3 == meltPtr_w ? _mask_ram_1_T : mask_ram_3_1; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_2_T = &io_inputBus_bits_mask_2; // @[WDB.scala 172:69]
  wire  _GEN_78 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_2 : mask_ram_0_2; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_79 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_2 : mask_ram_1_2; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_80 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_2 : mask_ram_2_2; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_81 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_2 : mask_ram_3_2; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_82 = 2'h0 == meltPtr_w ? _mask_ram_2_T : mask_ram_0_2; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_83 = 2'h1 == meltPtr_w ? _mask_ram_2_T : mask_ram_1_2; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_84 = 2'h2 == meltPtr_w ? _mask_ram_2_T : mask_ram_2_2; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_85 = 2'h3 == meltPtr_w ? _mask_ram_2_T : mask_ram_3_2; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_3_T = &io_inputBus_bits_mask_3; // @[WDB.scala 172:69]
  wire  _GEN_98 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_3 : mask_ram_0_3; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_99 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_3 : mask_ram_1_3; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_100 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_3 : mask_ram_2_3; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_101 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_3 : mask_ram_3_3; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_102 = 2'h0 == meltPtr_w ? _mask_ram_3_T : mask_ram_0_3; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_103 = 2'h1 == meltPtr_w ? _mask_ram_3_T : mask_ram_1_3; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_104 = 2'h2 == meltPtr_w ? _mask_ram_3_T : mask_ram_2_3; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_105 = 2'h3 == meltPtr_w ? _mask_ram_3_T : mask_ram_3_3; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_4_T = &io_inputBus_bits_mask_4; // @[WDB.scala 172:69]
  wire  _GEN_118 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_4 : mask_ram_0_4; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_119 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_4 : mask_ram_1_4; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_120 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_4 : mask_ram_2_4; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_121 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_4 : mask_ram_3_4; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_122 = 2'h0 == meltPtr_w ? _mask_ram_4_T : mask_ram_0_4; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_123 = 2'h1 == meltPtr_w ? _mask_ram_4_T : mask_ram_1_4; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_124 = 2'h2 == meltPtr_w ? _mask_ram_4_T : mask_ram_2_4; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_125 = 2'h3 == meltPtr_w ? _mask_ram_4_T : mask_ram_3_4; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_5_T = &io_inputBus_bits_mask_5; // @[WDB.scala 172:69]
  wire  _GEN_138 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_5 : mask_ram_0_5; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_139 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_5 : mask_ram_1_5; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_140 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_5 : mask_ram_2_5; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_141 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_5 : mask_ram_3_5; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_142 = 2'h0 == meltPtr_w ? _mask_ram_5_T : mask_ram_0_5; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_143 = 2'h1 == meltPtr_w ? _mask_ram_5_T : mask_ram_1_5; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_144 = 2'h2 == meltPtr_w ? _mask_ram_5_T : mask_ram_2_5; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_145 = 2'h3 == meltPtr_w ? _mask_ram_5_T : mask_ram_3_5; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_6_T = &io_inputBus_bits_mask_6; // @[WDB.scala 172:69]
  wire  _GEN_158 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_6 : mask_ram_0_6; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_159 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_6 : mask_ram_1_6; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_160 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_6 : mask_ram_2_6; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_161 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_6 : mask_ram_3_6; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_162 = 2'h0 == meltPtr_w ? _mask_ram_6_T : mask_ram_0_6; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_163 = 2'h1 == meltPtr_w ? _mask_ram_6_T : mask_ram_1_6; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_164 = 2'h2 == meltPtr_w ? _mask_ram_6_T : mask_ram_2_6; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_165 = 2'h3 == meltPtr_w ? _mask_ram_6_T : mask_ram_3_6; // @[WDB.scala 104:25 174:{35,35}]
  wire  _mask_ram_7_T = &io_inputBus_bits_mask_7; // @[WDB.scala 172:69]
  wire  _GEN_178 = 2'h0 == enqPtr_w ? &io_inputBus_bits_mask_7 : mask_ram_0_7; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_179 = 2'h1 == enqPtr_w ? &io_inputBus_bits_mask_7 : mask_ram_1_7; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_180 = 2'h2 == enqPtr_w ? &io_inputBus_bits_mask_7 : mask_ram_2_7; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_181 = 2'h3 == enqPtr_w ? &io_inputBus_bits_mask_7 : mask_ram_3_7; // @[WDB.scala 104:25 172:{34,34}]
  wire  _GEN_182 = 2'h0 == meltPtr_w ? _mask_ram_7_T : mask_ram_0_7; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_183 = 2'h1 == meltPtr_w ? _mask_ram_7_T : mask_ram_1_7; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_184 = 2'h2 == meltPtr_w ? _mask_ram_7_T : mask_ram_2_7; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_185 = 2'h3 == meltPtr_w ? _mask_ram_7_T : mask_ram_3_7; // @[WDB.scala 104:25 174:{35,35}]
  wire  _GEN_635 = 2'h1 == deqPtr_w ? mask_ram_1_0 : mask_ram_0_0; // @[WDB.scala 197:{26,26}]
  wire  _GEN_636 = 2'h2 == deqPtr_w ? mask_ram_2_0 : _GEN_635; // @[WDB.scala 197:{26,26}]
  wire  _GEN_639 = 2'h1 == deqPtr_w ? mask_ram_1_1 : mask_ram_0_1; // @[WDB.scala 197:{26,26}]
  wire  _GEN_640 = 2'h2 == deqPtr_w ? mask_ram_2_1 : _GEN_639; // @[WDB.scala 197:{26,26}]
  wire  _GEN_643 = 2'h1 == deqPtr_w ? mask_ram_1_2 : mask_ram_0_2; // @[WDB.scala 197:{26,26}]
  wire  _GEN_644 = 2'h2 == deqPtr_w ? mask_ram_2_2 : _GEN_643; // @[WDB.scala 197:{26,26}]
  wire  _GEN_647 = 2'h1 == deqPtr_w ? mask_ram_1_3 : mask_ram_0_3; // @[WDB.scala 197:{26,26}]
  wire  _GEN_648 = 2'h2 == deqPtr_w ? mask_ram_2_3 : _GEN_647; // @[WDB.scala 197:{26,26}]
  wire  _GEN_651 = 2'h1 == deqPtr_w ? mask_ram_1_4 : mask_ram_0_4; // @[WDB.scala 197:{26,26}]
  wire  _GEN_652 = 2'h2 == deqPtr_w ? mask_ram_2_4 : _GEN_651; // @[WDB.scala 197:{26,26}]
  wire  _GEN_655 = 2'h1 == deqPtr_w ? mask_ram_1_5 : mask_ram_0_5; // @[WDB.scala 197:{26,26}]
  wire  _GEN_656 = 2'h2 == deqPtr_w ? mask_ram_2_5 : _GEN_655; // @[WDB.scala 197:{26,26}]
  wire  _GEN_659 = 2'h1 == deqPtr_w ? mask_ram_1_6 : mask_ram_0_6; // @[WDB.scala 197:{26,26}]
  wire  _GEN_660 = 2'h2 == deqPtr_w ? mask_ram_2_6 : _GEN_659; // @[WDB.scala 197:{26,26}]
  wire  _GEN_663 = 2'h1 == deqPtr_w ? mask_ram_1_7 : mask_ram_0_7; // @[WDB.scala 197:{26,26}]
  wire  _GEN_664 = 2'h2 == deqPtr_w ? mask_ram_2_7 : _GEN_663; // @[WDB.scala 197:{26,26}]
  wire [31:0] _GEN_667 = 2'h1 == deqPtr_w ? addr_ram_1 : addr_ram_0; // @[WDB.scala 198:{26,26}]
  wire [31:0] _GEN_668 = 2'h2 == deqPtr_w ? addr_ram_2 : _GEN_667; // @[WDB.scala 198:{26,26}]
  wire [7:0] _GEN_671 = 2'h1 == deqPtr_w ? data_ram_1_0_0 : data_ram_0_0_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_672 = 2'h2 == deqPtr_w ? data_ram_2_0_0 : _GEN_671; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_675 = 2'h1 == deqPtr_w ? data_ram_1_0_1 : data_ram_0_0_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_676 = 2'h2 == deqPtr_w ? data_ram_2_0_1 : _GEN_675; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_679 = 2'h1 == deqPtr_w ? data_ram_1_0_2 : data_ram_0_0_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_680 = 2'h2 == deqPtr_w ? data_ram_2_0_2 : _GEN_679; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_683 = 2'h1 == deqPtr_w ? data_ram_1_0_3 : data_ram_0_0_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_684 = 2'h2 == deqPtr_w ? data_ram_2_0_3 : _GEN_683; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_687 = 2'h1 == deqPtr_w ? data_ram_1_1_0 : data_ram_0_1_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_688 = 2'h2 == deqPtr_w ? data_ram_2_1_0 : _GEN_687; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_691 = 2'h1 == deqPtr_w ? data_ram_1_1_1 : data_ram_0_1_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_692 = 2'h2 == deqPtr_w ? data_ram_2_1_1 : _GEN_691; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_695 = 2'h1 == deqPtr_w ? data_ram_1_1_2 : data_ram_0_1_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_696 = 2'h2 == deqPtr_w ? data_ram_2_1_2 : _GEN_695; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_699 = 2'h1 == deqPtr_w ? data_ram_1_1_3 : data_ram_0_1_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_700 = 2'h2 == deqPtr_w ? data_ram_2_1_3 : _GEN_699; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_703 = 2'h1 == deqPtr_w ? data_ram_1_2_0 : data_ram_0_2_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_704 = 2'h2 == deqPtr_w ? data_ram_2_2_0 : _GEN_703; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_707 = 2'h1 == deqPtr_w ? data_ram_1_2_1 : data_ram_0_2_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_708 = 2'h2 == deqPtr_w ? data_ram_2_2_1 : _GEN_707; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_711 = 2'h1 == deqPtr_w ? data_ram_1_2_2 : data_ram_0_2_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_712 = 2'h2 == deqPtr_w ? data_ram_2_2_2 : _GEN_711; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_715 = 2'h1 == deqPtr_w ? data_ram_1_2_3 : data_ram_0_2_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_716 = 2'h2 == deqPtr_w ? data_ram_2_2_3 : _GEN_715; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_719 = 2'h1 == deqPtr_w ? data_ram_1_3_0 : data_ram_0_3_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_720 = 2'h2 == deqPtr_w ? data_ram_2_3_0 : _GEN_719; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_723 = 2'h1 == deqPtr_w ? data_ram_1_3_1 : data_ram_0_3_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_724 = 2'h2 == deqPtr_w ? data_ram_2_3_1 : _GEN_723; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_727 = 2'h1 == deqPtr_w ? data_ram_1_3_2 : data_ram_0_3_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_728 = 2'h2 == deqPtr_w ? data_ram_2_3_2 : _GEN_727; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_731 = 2'h1 == deqPtr_w ? data_ram_1_3_3 : data_ram_0_3_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_732 = 2'h2 == deqPtr_w ? data_ram_2_3_3 : _GEN_731; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_735 = 2'h1 == deqPtr_w ? data_ram_1_4_0 : data_ram_0_4_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_736 = 2'h2 == deqPtr_w ? data_ram_2_4_0 : _GEN_735; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_739 = 2'h1 == deqPtr_w ? data_ram_1_4_1 : data_ram_0_4_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_740 = 2'h2 == deqPtr_w ? data_ram_2_4_1 : _GEN_739; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_743 = 2'h1 == deqPtr_w ? data_ram_1_4_2 : data_ram_0_4_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_744 = 2'h2 == deqPtr_w ? data_ram_2_4_2 : _GEN_743; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_747 = 2'h1 == deqPtr_w ? data_ram_1_4_3 : data_ram_0_4_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_748 = 2'h2 == deqPtr_w ? data_ram_2_4_3 : _GEN_747; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_751 = 2'h1 == deqPtr_w ? data_ram_1_5_0 : data_ram_0_5_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_752 = 2'h2 == deqPtr_w ? data_ram_2_5_0 : _GEN_751; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_755 = 2'h1 == deqPtr_w ? data_ram_1_5_1 : data_ram_0_5_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_756 = 2'h2 == deqPtr_w ? data_ram_2_5_1 : _GEN_755; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_759 = 2'h1 == deqPtr_w ? data_ram_1_5_2 : data_ram_0_5_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_760 = 2'h2 == deqPtr_w ? data_ram_2_5_2 : _GEN_759; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_763 = 2'h1 == deqPtr_w ? data_ram_1_5_3 : data_ram_0_5_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_764 = 2'h2 == deqPtr_w ? data_ram_2_5_3 : _GEN_763; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_767 = 2'h1 == deqPtr_w ? data_ram_1_6_0 : data_ram_0_6_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_768 = 2'h2 == deqPtr_w ? data_ram_2_6_0 : _GEN_767; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_771 = 2'h1 == deqPtr_w ? data_ram_1_6_1 : data_ram_0_6_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_772 = 2'h2 == deqPtr_w ? data_ram_2_6_1 : _GEN_771; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_775 = 2'h1 == deqPtr_w ? data_ram_1_6_2 : data_ram_0_6_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_776 = 2'h2 == deqPtr_w ? data_ram_2_6_2 : _GEN_775; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_779 = 2'h1 == deqPtr_w ? data_ram_1_6_3 : data_ram_0_6_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_780 = 2'h2 == deqPtr_w ? data_ram_2_6_3 : _GEN_779; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_783 = 2'h1 == deqPtr_w ? data_ram_1_7_0 : data_ram_0_7_0; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_784 = 2'h2 == deqPtr_w ? data_ram_2_7_0 : _GEN_783; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_787 = 2'h1 == deqPtr_w ? data_ram_1_7_1 : data_ram_0_7_1; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_788 = 2'h2 == deqPtr_w ? data_ram_2_7_1 : _GEN_787; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_791 = 2'h1 == deqPtr_w ? data_ram_1_7_2 : data_ram_0_7_2; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_792 = 2'h2 == deqPtr_w ? data_ram_2_7_2 : _GEN_791; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_795 = 2'h1 == deqPtr_w ? data_ram_1_7_3 : data_ram_0_7_3; // @[WDB.scala 199:{26,26}]
  wire [7:0] _GEN_796 = 2'h2 == deqPtr_w ? data_ram_2_7_3 : _GEN_795; // @[WDB.scala 199:{26,26}]
  wire [1:0] _GEN_799 = 2'h1 == deqPtr_w ? instrId_ram_1 : instrId_ram_0; // @[WDB.scala 200:{29,29}]
  wire [1:0] _GEN_800 = 2'h2 == deqPtr_w ? instrId_ram_2 : _GEN_799; // @[WDB.scala 200:{29,29}]
  wire  full = _almFull_T_9 == 3'h4; // @[WDB.scala 203:40]
  wire [3:0] _unfrozenCount_T_1 = {entryFrozen_0,entryFrozen_1,entryFrozen_2,entryFrozen_3}; // @[Cat.scala 31:58]
  wire [3:0] _unfrozenCount_T_2 = _almFull_T ^ _unfrozenCount_T_1; // @[WDB.scala 207:47]
  wire [1:0] _unfrozenCount_T_7 = _unfrozenCount_T_2[0] + _unfrozenCount_T_2[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _unfrozenCount_T_9 = _unfrozenCount_T_2[2] + _unfrozenCount_T_2[3]; // @[Bitwise.scala 48:55]
  wire [2:0] unfrozenCount = _unfrozenCount_T_7 + _unfrozenCount_T_9; // @[Bitwise.scala 48:55]
  wire  empty = unfrozenCount == 3'h0; // @[WDB.scala 208:29]
  wire [2:0] _io_wdbAlmostFull_T_1 = 3'h4 - 3'h2; // @[WDB.scala 210:59]
  WdbEnqPtrGen enqPtr_w_Gen ( // @[WDB.scala 53:21]
    .io_entryValidList_0(enqPtr_w_Gen_io_entryValidList_0),
    .io_entryValidList_1(enqPtr_w_Gen_io_entryValidList_1),
    .io_entryValidList_2(enqPtr_w_Gen_io_entryValidList_2),
    .io_entryValidList_3(enqPtr_w_Gen_io_entryValidList_3),
    .io_enqPtr_cs(enqPtr_w_Gen_io_enqPtr_cs),
    .io_enqPtr_ns(enqPtr_w_Gen_io_enqPtr_ns)
  );
  WdbDeqPtrGen deqPtr_w_Gen ( // @[WDB.scala 89:21]
    .io_entryValidList_0(deqPtr_w_Gen_io_entryValidList_0),
    .io_entryValidList_1(deqPtr_w_Gen_io_entryValidList_1),
    .io_entryValidList_2(deqPtr_w_Gen_io_entryValidList_2),
    .io_entryValidList_3(deqPtr_w_Gen_io_entryValidList_3),
    .io_entryFrozenList_0(deqPtr_w_Gen_io_entryFrozenList_0),
    .io_entryFrozenList_1(deqPtr_w_Gen_io_entryFrozenList_1),
    .io_entryFrozenList_2(deqPtr_w_Gen_io_entryFrozenList_2),
    .io_entryFrozenList_3(deqPtr_w_Gen_io_entryFrozenList_3),
    .io_deqPtr_cs(deqPtr_w_Gen_io_deqPtr_cs),
    .io_deqPtr_ns(deqPtr_w_Gen_io_deqPtr_ns)
  );
  assign io_inputBus_ready = ~full; // @[WDB.scala 204:24]
  assign io_outputBus_valid = ~empty; // @[WDB.scala 209:25]
  assign io_outputBus_bits_mask_0 = 2'h3 == deqPtr_w ? mask_ram_3_0 : _GEN_636; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_1 = 2'h3 == deqPtr_w ? mask_ram_3_1 : _GEN_640; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_2 = 2'h3 == deqPtr_w ? mask_ram_3_2 : _GEN_644; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_3 = 2'h3 == deqPtr_w ? mask_ram_3_3 : _GEN_648; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_4 = 2'h3 == deqPtr_w ? mask_ram_3_4 : _GEN_652; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_5 = 2'h3 == deqPtr_w ? mask_ram_3_5 : _GEN_656; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_6 = 2'h3 == deqPtr_w ? mask_ram_3_6 : _GEN_660; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_mask_7 = 2'h3 == deqPtr_w ? mask_ram_3_7 : _GEN_664; // @[WDB.scala 197:{26,26}]
  assign io_outputBus_bits_addr = 2'h3 == deqPtr_w ? addr_ram_3 : _GEN_668; // @[WDB.scala 198:{26,26}]
  assign io_outputBus_bits_data_0_0 = 2'h3 == deqPtr_w ? data_ram_3_0_0 : _GEN_672; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_0_1 = 2'h3 == deqPtr_w ? data_ram_3_0_1 : _GEN_676; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_0_2 = 2'h3 == deqPtr_w ? data_ram_3_0_2 : _GEN_680; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_0_3 = 2'h3 == deqPtr_w ? data_ram_3_0_3 : _GEN_684; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_1_0 = 2'h3 == deqPtr_w ? data_ram_3_1_0 : _GEN_688; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_1_1 = 2'h3 == deqPtr_w ? data_ram_3_1_1 : _GEN_692; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_1_2 = 2'h3 == deqPtr_w ? data_ram_3_1_2 : _GEN_696; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_1_3 = 2'h3 == deqPtr_w ? data_ram_3_1_3 : _GEN_700; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_2_0 = 2'h3 == deqPtr_w ? data_ram_3_2_0 : _GEN_704; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_2_1 = 2'h3 == deqPtr_w ? data_ram_3_2_1 : _GEN_708; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_2_2 = 2'h3 == deqPtr_w ? data_ram_3_2_2 : _GEN_712; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_2_3 = 2'h3 == deqPtr_w ? data_ram_3_2_3 : _GEN_716; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_3_0 = 2'h3 == deqPtr_w ? data_ram_3_3_0 : _GEN_720; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_3_1 = 2'h3 == deqPtr_w ? data_ram_3_3_1 : _GEN_724; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_3_2 = 2'h3 == deqPtr_w ? data_ram_3_3_2 : _GEN_728; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_3_3 = 2'h3 == deqPtr_w ? data_ram_3_3_3 : _GEN_732; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_4_0 = 2'h3 == deqPtr_w ? data_ram_3_4_0 : _GEN_736; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_4_1 = 2'h3 == deqPtr_w ? data_ram_3_4_1 : _GEN_740; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_4_2 = 2'h3 == deqPtr_w ? data_ram_3_4_2 : _GEN_744; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_4_3 = 2'h3 == deqPtr_w ? data_ram_3_4_3 : _GEN_748; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_5_0 = 2'h3 == deqPtr_w ? data_ram_3_5_0 : _GEN_752; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_5_1 = 2'h3 == deqPtr_w ? data_ram_3_5_1 : _GEN_756; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_5_2 = 2'h3 == deqPtr_w ? data_ram_3_5_2 : _GEN_760; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_5_3 = 2'h3 == deqPtr_w ? data_ram_3_5_3 : _GEN_764; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_6_0 = 2'h3 == deqPtr_w ? data_ram_3_6_0 : _GEN_768; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_6_1 = 2'h3 == deqPtr_w ? data_ram_3_6_1 : _GEN_772; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_6_2 = 2'h3 == deqPtr_w ? data_ram_3_6_2 : _GEN_776; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_6_3 = 2'h3 == deqPtr_w ? data_ram_3_6_3 : _GEN_780; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_7_0 = 2'h3 == deqPtr_w ? data_ram_3_7_0 : _GEN_784; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_7_1 = 2'h3 == deqPtr_w ? data_ram_3_7_1 : _GEN_788; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_7_2 = 2'h3 == deqPtr_w ? data_ram_3_7_2 : _GEN_792; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_data_7_3 = 2'h3 == deqPtr_w ? data_ram_3_7_3 : _GEN_796; // @[WDB.scala 199:{26,26}]
  assign io_outputBus_bits_instrId = 2'h3 == deqPtr_w ? instrId_ram_3 : _GEN_800; // @[WDB.scala 200:{29,29}]
  assign io_wdbAlmostFull = unfrozenCount == _io_wdbAlmostFull_T_1; // @[WDB.scala 210:37]
  assign enqPtr_w_Gen_io_entryValidList_0 = entryValid_0; // @[WDB.scala 54:27]
  assign enqPtr_w_Gen_io_entryValidList_1 = entryValid_1; // @[WDB.scala 54:27]
  assign enqPtr_w_Gen_io_entryValidList_2 = entryValid_2; // @[WDB.scala 54:27]
  assign enqPtr_w_Gen_io_entryValidList_3 = entryValid_3; // @[WDB.scala 54:27]
  assign enqPtr_w_Gen_io_enqPtr_cs = enqPtr; // @[WDB.scala 55:22]
  assign deqPtr_w_Gen_io_entryValidList_0 = entryValid_0; // @[WDB.scala 90:27]
  assign deqPtr_w_Gen_io_entryValidList_1 = entryValid_1; // @[WDB.scala 90:27]
  assign deqPtr_w_Gen_io_entryValidList_2 = entryValid_2; // @[WDB.scala 90:27]
  assign deqPtr_w_Gen_io_entryValidList_3 = entryValid_3; // @[WDB.scala 90:27]
  assign deqPtr_w_Gen_io_entryFrozenList_0 = entryFrozen_0; // @[WDB.scala 91:28]
  assign deqPtr_w_Gen_io_entryFrozenList_1 = entryFrozen_1; // @[WDB.scala 91:28]
  assign deqPtr_w_Gen_io_entryFrozenList_2 = entryFrozen_2; // @[WDB.scala 91:28]
  assign deqPtr_w_Gen_io_entryFrozenList_3 = entryFrozen_3; // @[WDB.scala 91:28]
  assign deqPtr_w_Gen_io_deqPtr_cs = deqPtr; // @[WDB.scala 92:22]
  always @(posedge clock) begin
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_0 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_0 <= _GEN_38;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_0 <= _GEN_42;
      end else begin
        mask_ram_0_0 <= _GEN_38;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_1 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_1 <= _GEN_58;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_1 <= _GEN_62;
      end else begin
        mask_ram_0_1 <= _GEN_58;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_2 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_2 <= _GEN_78;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_2 <= _GEN_82;
      end else begin
        mask_ram_0_2 <= _GEN_78;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_3 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_3 <= _GEN_98;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_3 <= _GEN_102;
      end else begin
        mask_ram_0_3 <= _GEN_98;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_4 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_4 <= _GEN_118;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_4 <= _GEN_122;
      end else begin
        mask_ram_0_4 <= _GEN_118;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_5 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_5 <= _GEN_138;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_5 <= _GEN_142;
      end else begin
        mask_ram_0_5 <= _GEN_138;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_6 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_6 <= _GEN_158;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_6 <= _GEN_162;
      end else begin
        mask_ram_0_6 <= _GEN_158;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_0_7 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_0_7 <= _GEN_178;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_0_7 <= _GEN_182;
      end else begin
        mask_ram_0_7 <= _GEN_178;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_0 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_0 <= _GEN_39;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_0 <= _GEN_43;
      end else begin
        mask_ram_1_0 <= _GEN_39;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_1 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_1 <= _GEN_59;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_1 <= _GEN_63;
      end else begin
        mask_ram_1_1 <= _GEN_59;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_2 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_2 <= _GEN_79;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_2 <= _GEN_83;
      end else begin
        mask_ram_1_2 <= _GEN_79;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_3 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_3 <= _GEN_99;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_3 <= _GEN_103;
      end else begin
        mask_ram_1_3 <= _GEN_99;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_4 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_4 <= _GEN_119;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_4 <= _GEN_123;
      end else begin
        mask_ram_1_4 <= _GEN_119;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_5 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_5 <= _GEN_139;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_5 <= _GEN_143;
      end else begin
        mask_ram_1_5 <= _GEN_139;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_6 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_6 <= _GEN_159;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_6 <= _GEN_163;
      end else begin
        mask_ram_1_6 <= _GEN_159;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_1_7 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_1_7 <= _GEN_179;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_1_7 <= _GEN_183;
      end else begin
        mask_ram_1_7 <= _GEN_179;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_0 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_0 <= _GEN_40;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_0 <= _GEN_44;
      end else begin
        mask_ram_2_0 <= _GEN_40;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_1 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_1 <= _GEN_60;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_1 <= _GEN_64;
      end else begin
        mask_ram_2_1 <= _GEN_60;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_2 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_2 <= _GEN_80;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_2 <= _GEN_84;
      end else begin
        mask_ram_2_2 <= _GEN_80;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_3 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_3 <= _GEN_100;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_3 <= _GEN_104;
      end else begin
        mask_ram_2_3 <= _GEN_100;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_4 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_4 <= _GEN_120;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_4 <= _GEN_124;
      end else begin
        mask_ram_2_4 <= _GEN_120;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_5 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_5 <= _GEN_140;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_5 <= _GEN_144;
      end else begin
        mask_ram_2_5 <= _GEN_140;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_6 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_6 <= _GEN_160;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_6 <= _GEN_164;
      end else begin
        mask_ram_2_6 <= _GEN_160;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_2_7 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_2_7 <= _GEN_180;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_2_7 <= _GEN_184;
      end else begin
        mask_ram_2_7 <= _GEN_180;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_0 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_0 <= _GEN_41;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_0 <= _GEN_45;
      end else begin
        mask_ram_3_0 <= _GEN_41;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_1 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_1 <= _GEN_61;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_1 <= _GEN_65;
      end else begin
        mask_ram_3_1 <= _GEN_61;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_2 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_2 <= _GEN_81;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_2 <= _GEN_85;
      end else begin
        mask_ram_3_2 <= _GEN_81;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_3 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_3 <= _GEN_101;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_3 <= _GEN_105;
      end else begin
        mask_ram_3_3 <= _GEN_101;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_4 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_4 <= _GEN_121;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_4 <= _GEN_125;
      end else begin
        mask_ram_3_4 <= _GEN_121;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_5 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_5 <= _GEN_141;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_5 <= _GEN_145;
      end else begin
        mask_ram_3_5 <= _GEN_141;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_6 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_6 <= _GEN_161;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_6 <= _GEN_165;
      end else begin
        mask_ram_3_6 <= _GEN_161;
      end
    end
    if (reset) begin // @[WDB.scala 104:25]
      mask_ram_3_7 <= 1'h0; // @[WDB.scala 104:25]
    end else if (doEnq) begin // @[WDB.scala 169:15]
      if (io_inputBus_bits_subWordMissReq) begin // @[WDB.scala 171:27]
        mask_ram_3_7 <= _GEN_181;
      end else if (io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 173:33]
        mask_ram_3_7 <= _GEN_185;
      end else begin
        mask_ram_3_7 <= _GEN_181;
      end
    end
    if (reset) begin // @[WDB.scala 105:25]
      addr_ram_0 <= 32'h0; // @[WDB.scala 105:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (_T_15) begin // @[WDB.scala 191:27]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 192:26]
          addr_ram_0 <= io_inputBus_bits_addr; // @[WDB.scala 192:26]
        end
      end
    end
    if (reset) begin // @[WDB.scala 105:25]
      addr_ram_1 <= 32'h0; // @[WDB.scala 105:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (_T_15) begin // @[WDB.scala 191:27]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 192:26]
          addr_ram_1 <= io_inputBus_bits_addr; // @[WDB.scala 192:26]
        end
      end
    end
    if (reset) begin // @[WDB.scala 105:25]
      addr_ram_2 <= 32'h0; // @[WDB.scala 105:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (_T_15) begin // @[WDB.scala 191:27]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 192:26]
          addr_ram_2 <= io_inputBus_bits_addr; // @[WDB.scala 192:26]
        end
      end
    end
    if (reset) begin // @[WDB.scala 105:25]
      addr_ram_3 <= 32'h0; // @[WDB.scala 105:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (_T_15) begin // @[WDB.scala 191:27]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 192:26]
          addr_ram_3 <= io_inputBus_bits_addr; // @[WDB.scala 192:26]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_0_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_0_0 <= io_inputBus_bits_data_0_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_0_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_0_1 <= io_inputBus_bits_data_0_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_0_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_0_2 <= io_inputBus_bits_data_0_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_0_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_0_3 <= io_inputBus_bits_data_0_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_1_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_1_0 <= io_inputBus_bits_data_1_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_1_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_1_1 <= io_inputBus_bits_data_1_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_1_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_1_2 <= io_inputBus_bits_data_1_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_1_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_1_3 <= io_inputBus_bits_data_1_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_2_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_2_0 <= io_inputBus_bits_data_2_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_2_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_2_1 <= io_inputBus_bits_data_2_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_2_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_2_2 <= io_inputBus_bits_data_2_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_2_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_2_3 <= io_inputBus_bits_data_2_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_3_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_3_0 <= io_inputBus_bits_data_3_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_3_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_3_1 <= io_inputBus_bits_data_3_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_3_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_3_2 <= io_inputBus_bits_data_3_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_3_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_3_3 <= io_inputBus_bits_data_3_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_4_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_4_0 <= io_inputBus_bits_data_4_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_4_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_4_1 <= io_inputBus_bits_data_4_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_4_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_4_2 <= io_inputBus_bits_data_4_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_4_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_4_3 <= io_inputBus_bits_data_4_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_5_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_5_0 <= io_inputBus_bits_data_5_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_5_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_5_1 <= io_inputBus_bits_data_5_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_5_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_5_2 <= io_inputBus_bits_data_5_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_5_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_5_3 <= io_inputBus_bits_data_5_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_6_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_6_0 <= io_inputBus_bits_data_6_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_6_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_6_1 <= io_inputBus_bits_data_6_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_6_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_6_2 <= io_inputBus_bits_data_6_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_6_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_6_3 <= io_inputBus_bits_data_6_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_7_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[0]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_7_0 <= io_inputBus_bits_data_7_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_7_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[1]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_7_1 <= io_inputBus_bits_data_7_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_7_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[2]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_7_2 <= io_inputBus_bits_data_7_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_0_7_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[3]) begin // @[WDB.scala 185:49]
        if (2'h0 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_0_7_3 <= io_inputBus_bits_data_7_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_0_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_0_0 <= io_inputBus_bits_data_0_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_0_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_0_1 <= io_inputBus_bits_data_0_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_0_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_0_2 <= io_inputBus_bits_data_0_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_0_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_0_3 <= io_inputBus_bits_data_0_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_1_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_1_0 <= io_inputBus_bits_data_1_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_1_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_1_1 <= io_inputBus_bits_data_1_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_1_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_1_2 <= io_inputBus_bits_data_1_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_1_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_1_3 <= io_inputBus_bits_data_1_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_2_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_2_0 <= io_inputBus_bits_data_2_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_2_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_2_1 <= io_inputBus_bits_data_2_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_2_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_2_2 <= io_inputBus_bits_data_2_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_2_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_2_3 <= io_inputBus_bits_data_2_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_3_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_3_0 <= io_inputBus_bits_data_3_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_3_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_3_1 <= io_inputBus_bits_data_3_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_3_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_3_2 <= io_inputBus_bits_data_3_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_3_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_3_3 <= io_inputBus_bits_data_3_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_4_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_4_0 <= io_inputBus_bits_data_4_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_4_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_4_1 <= io_inputBus_bits_data_4_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_4_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_4_2 <= io_inputBus_bits_data_4_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_4_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_4_3 <= io_inputBus_bits_data_4_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_5_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_5_0 <= io_inputBus_bits_data_5_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_5_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_5_1 <= io_inputBus_bits_data_5_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_5_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_5_2 <= io_inputBus_bits_data_5_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_5_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_5_3 <= io_inputBus_bits_data_5_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_6_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_6_0 <= io_inputBus_bits_data_6_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_6_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_6_1 <= io_inputBus_bits_data_6_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_6_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_6_2 <= io_inputBus_bits_data_6_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_6_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_6_3 <= io_inputBus_bits_data_6_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_7_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[0]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_7_0 <= io_inputBus_bits_data_7_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_7_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[1]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_7_1 <= io_inputBus_bits_data_7_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_7_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[2]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_7_2 <= io_inputBus_bits_data_7_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_1_7_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[3]) begin // @[WDB.scala 185:49]
        if (2'h1 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_1_7_3 <= io_inputBus_bits_data_7_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_0_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_0_0 <= io_inputBus_bits_data_0_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_0_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_0_1 <= io_inputBus_bits_data_0_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_0_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_0_2 <= io_inputBus_bits_data_0_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_0_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_0_3 <= io_inputBus_bits_data_0_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_1_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_1_0 <= io_inputBus_bits_data_1_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_1_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_1_1 <= io_inputBus_bits_data_1_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_1_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_1_2 <= io_inputBus_bits_data_1_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_1_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_1_3 <= io_inputBus_bits_data_1_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_2_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_2_0 <= io_inputBus_bits_data_2_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_2_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_2_1 <= io_inputBus_bits_data_2_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_2_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_2_2 <= io_inputBus_bits_data_2_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_2_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_2_3 <= io_inputBus_bits_data_2_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_3_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_3_0 <= io_inputBus_bits_data_3_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_3_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_3_1 <= io_inputBus_bits_data_3_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_3_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_3_2 <= io_inputBus_bits_data_3_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_3_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_3_3 <= io_inputBus_bits_data_3_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_4_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_4_0 <= io_inputBus_bits_data_4_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_4_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_4_1 <= io_inputBus_bits_data_4_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_4_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_4_2 <= io_inputBus_bits_data_4_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_4_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_4_3 <= io_inputBus_bits_data_4_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_5_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_5_0 <= io_inputBus_bits_data_5_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_5_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_5_1 <= io_inputBus_bits_data_5_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_5_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_5_2 <= io_inputBus_bits_data_5_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_5_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_5_3 <= io_inputBus_bits_data_5_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_6_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_6_0 <= io_inputBus_bits_data_6_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_6_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_6_1 <= io_inputBus_bits_data_6_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_6_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_6_2 <= io_inputBus_bits_data_6_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_6_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_6_3 <= io_inputBus_bits_data_6_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_7_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[0]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_7_0 <= io_inputBus_bits_data_7_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_7_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[1]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_7_1 <= io_inputBus_bits_data_7_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_7_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[2]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_7_2 <= io_inputBus_bits_data_7_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_2_7_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[3]) begin // @[WDB.scala 185:49]
        if (2'h2 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_2_7_3 <= io_inputBus_bits_data_7_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_0_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_0_0 <= io_inputBus_bits_data_0_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_0_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_0_1 <= io_inputBus_bits_data_0_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_0_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_0_2 <= io_inputBus_bits_data_0_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_0_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_0[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_0_3 <= io_inputBus_bits_data_0_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_1_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_1_0 <= io_inputBus_bits_data_1_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_1_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_1_1 <= io_inputBus_bits_data_1_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_1_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_1_2 <= io_inputBus_bits_data_1_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_1_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_1[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_1_3 <= io_inputBus_bits_data_1_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_2_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_2_0 <= io_inputBus_bits_data_2_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_2_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_2_1 <= io_inputBus_bits_data_2_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_2_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_2_2 <= io_inputBus_bits_data_2_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_2_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_2[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_2_3 <= io_inputBus_bits_data_2_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_3_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_3_0 <= io_inputBus_bits_data_3_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_3_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_3_1 <= io_inputBus_bits_data_3_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_3_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_3_2 <= io_inputBus_bits_data_3_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_3_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_3[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_3_3 <= io_inputBus_bits_data_3_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_4_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_4_0 <= io_inputBus_bits_data_4_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_4_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_4_1 <= io_inputBus_bits_data_4_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_4_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_4_2 <= io_inputBus_bits_data_4_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_4_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_4[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_4_3 <= io_inputBus_bits_data_4_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_5_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_5_0 <= io_inputBus_bits_data_5_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_5_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_5_1 <= io_inputBus_bits_data_5_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_5_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_5_2 <= io_inputBus_bits_data_5_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_5_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_5[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_5_3 <= io_inputBus_bits_data_5_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_6_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_6_0 <= io_inputBus_bits_data_6_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_6_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_6_1 <= io_inputBus_bits_data_6_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_6_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_6_2 <= io_inputBus_bits_data_6_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_6_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_6[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_6_3 <= io_inputBus_bits_data_6_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_7_0 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[0]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_7_0 <= io_inputBus_bits_data_7_0; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_7_1 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[1]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_7_1 <= io_inputBus_bits_data_7_1; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_7_2 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[2]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_7_2 <= io_inputBus_bits_data_7_2; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 106:25]
      data_ram_3_7_3 <= 8'h0; // @[WDB.scala 106:25]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (io_inputBus_bits_mask_7[3]) begin // @[WDB.scala 185:49]
        if (2'h3 == enqPtr_w) begin // @[WDB.scala 186:42]
          data_ram_3_7_3 <= io_inputBus_bits_data_7_3; // @[WDB.scala 186:42]
        end
      end
    end
    if (reset) begin // @[WDB.scala 109:28]
      instrId_ram_0 <= 2'h0; // @[WDB.scala 109:28]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (2'h0 == enqPtr_w) begin // @[WDB.scala 190:27]
        instrId_ram_0 <= io_inputBus_bits_instrId; // @[WDB.scala 190:27]
      end
    end
    if (reset) begin // @[WDB.scala 109:28]
      instrId_ram_1 <= 2'h0; // @[WDB.scala 109:28]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (2'h1 == enqPtr_w) begin // @[WDB.scala 190:27]
        instrId_ram_1 <= io_inputBus_bits_instrId; // @[WDB.scala 190:27]
      end
    end
    if (reset) begin // @[WDB.scala 109:28]
      instrId_ram_2 <= 2'h0; // @[WDB.scala 109:28]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (2'h2 == enqPtr_w) begin // @[WDB.scala 190:27]
        instrId_ram_2 <= io_inputBus_bits_instrId; // @[WDB.scala 190:27]
      end
    end
    if (reset) begin // @[WDB.scala 109:28]
      instrId_ram_3 <= 2'h0; // @[WDB.scala 109:28]
    end else if (doEnq) begin // @[WDB.scala 182:15]
      if (2'h3 == enqPtr_w) begin // @[WDB.scala 190:27]
        instrId_ram_3 <= io_inputBus_bits_instrId; // @[WDB.scala 190:27]
      end
    end
    if (reset) begin // @[WDB.scala 111:23]
      enqPtr <= 2'h0; // @[WDB.scala 111:23]
    end else if (doEnq & ~io_inputBus_bits_bankConflict) begin // @[WDB.scala 133:33]
      enqPtr <= enqPtr_w; // @[WDB.scala 134:12]
    end
    if (reset) begin // @[WDB.scala 112:23]
      deqPtr <= 2'h0; // @[WDB.scala 112:23]
    end else if (doDeq) begin // @[WDB.scala 138:15]
      deqPtr <= deqPtr_w; // @[WDB.scala 139:12]
    end
    if (reset) begin // @[WDB.scala 118:27]
      entryValid_0 <= 1'h0; // @[WDB.scala 118:27]
    end else if (2'h0 == deqPtr_w & doDeq) begin // @[WDB.scala 152:39]
      entryValid_0 <= 1'h0; // @[WDB.scala 154:21]
    end else if (_T_1) begin // @[WDB.scala 155:40]
      entryValid_0 <= _GEN_7;
    end
    if (reset) begin // @[WDB.scala 118:27]
      entryValid_1 <= 1'h0; // @[WDB.scala 118:27]
    end else if (2'h1 == deqPtr_w & doDeq) begin // @[WDB.scala 152:39]
      entryValid_1 <= 1'h0; // @[WDB.scala 154:21]
    end else if (_T_1) begin // @[WDB.scala 155:40]
      entryValid_1 <= _GEN_15;
    end
    if (reset) begin // @[WDB.scala 118:27]
      entryValid_2 <= 1'h0; // @[WDB.scala 118:27]
    end else if (2'h2 == deqPtr_w & doDeq) begin // @[WDB.scala 152:39]
      entryValid_2 <= 1'h0; // @[WDB.scala 154:21]
    end else if (_T_1) begin // @[WDB.scala 155:40]
      entryValid_2 <= _GEN_23;
    end
    if (reset) begin // @[WDB.scala 118:27]
      entryValid_3 <= 1'h0; // @[WDB.scala 118:27]
    end else if (2'h3 == deqPtr_w & doDeq) begin // @[WDB.scala 152:39]
      entryValid_3 <= 1'h0; // @[WDB.scala 154:21]
    end else if (_T_1) begin // @[WDB.scala 155:40]
      entryValid_3 <= _GEN_31;
    end
    if (reset) begin // @[WDB.scala 119:28]
      entryFrozen_0 <= 1'h0; // @[WDB.scala 119:28]
    end else if (!(2'h0 == deqPtr_w & doDeq)) begin // @[WDB.scala 152:39]
      if (_T_1) begin // @[WDB.scala 155:40]
        if (2'h0 == meltPtr_w & io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 162:51]
          entryFrozen_0 <= 1'h0; // @[WDB.scala 163:24]
        end else begin
          entryFrozen_0 <= _GEN_8;
        end
      end
    end
    if (reset) begin // @[WDB.scala 119:28]
      entryFrozen_1 <= 1'h0; // @[WDB.scala 119:28]
    end else if (!(2'h1 == deqPtr_w & doDeq)) begin // @[WDB.scala 152:39]
      if (_T_1) begin // @[WDB.scala 155:40]
        if (2'h1 == meltPtr_w & io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 162:51]
          entryFrozen_1 <= 1'h0; // @[WDB.scala 163:24]
        end else begin
          entryFrozen_1 <= _GEN_16;
        end
      end
    end
    if (reset) begin // @[WDB.scala 119:28]
      entryFrozen_2 <= 1'h0; // @[WDB.scala 119:28]
    end else if (!(2'h2 == deqPtr_w & doDeq)) begin // @[WDB.scala 152:39]
      if (_T_1) begin // @[WDB.scala 155:40]
        if (2'h2 == meltPtr_w & io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 162:51]
          entryFrozen_2 <= 1'h0; // @[WDB.scala 163:24]
        end else begin
          entryFrozen_2 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[WDB.scala 119:28]
      entryFrozen_3 <= 1'h0; // @[WDB.scala 119:28]
    end else if (!(2'h3 == deqPtr_w & doDeq)) begin // @[WDB.scala 152:39]
      if (_T_1) begin // @[WDB.scala 155:40]
        if (2'h3 == meltPtr_w & io_inputBus_bits_subWordMissRsp) begin // @[WDB.scala 162:51]
          entryFrozen_3 <= 1'h0; // @[WDB.scala 163:24]
        end else begin
          entryFrozen_3 <= _GEN_32;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(_T_11 == 3'h1 & io_inputBus_bits_subWordMissRsp | ~io_inputBus_bits_subWordMissRsp)) begin
          $fatal; // @[WDB.scala 146:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_11 == 3'h1 & io_inputBus_bits_subWordMissRsp | ~io_inputBus_bits_subWordMissRsp)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:146 assert((PopCount(Cat(meltMatch))===1.U && subWordMissRsp) || !subWordMissRsp)\n"
            ); // @[WDB.scala 146:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_18 & ~(_GEN_5 & io_inputBus_bits_subWordMissRsp | _T_15)) begin
          $fatal; // @[WDB.scala 148:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_18 & ~(_GEN_5 & io_inputBus_bits_subWordMissRsp | _T_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:148 assert((entryFrozen(meltPtr_w)===true.B && subWordMissRsp) || !subWordMissRsp)\n"
            ); // @[WDB.scala 148:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_0 == _mask_ram_0_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_0 == _mask_ram_0_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_1 == _mask_ram_1_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_1 == _mask_ram_1_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_2 == _mask_ram_2_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_2 == _mask_ram_2_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_3 == _mask_ram_3_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_3 == _mask_ram_3_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_4 == _mask_ram_4_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_4 == _mask_ram_4_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_5 == _mask_ram_5_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_5 == _mask_ram_5_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_6 == _mask_ram_6_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_6 == _mask_ram_6_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_7 == _mask_ram_7_T)
          ) begin
          $fatal; // @[WDB.scala 177:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doEnq & ~io_inputBus_bits_subWordMissReq & _T_15 & _T_18 & ~(|io_inputBus_bits_mask_7 == _mask_ram_7_T)
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WDB.scala:177 assert(io.inputBus.bits.mask(iofW).orR === io.inputBus.bits.mask(iofW).andR)\n"
            ); // @[WDB.scala 177:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mask_ram_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mask_ram_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mask_ram_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  mask_ram_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  mask_ram_0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  mask_ram_0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mask_ram_0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  mask_ram_0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mask_ram_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mask_ram_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  mask_ram_1_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  mask_ram_1_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  mask_ram_1_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  mask_ram_1_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  mask_ram_1_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  mask_ram_1_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  mask_ram_2_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  mask_ram_2_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  mask_ram_2_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  mask_ram_2_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mask_ram_2_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  mask_ram_2_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  mask_ram_2_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  mask_ram_2_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  mask_ram_3_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  mask_ram_3_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  mask_ram_3_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  mask_ram_3_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mask_ram_3_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  mask_ram_3_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  mask_ram_3_6 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  mask_ram_3_7 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  addr_ram_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  addr_ram_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  addr_ram_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  addr_ram_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  data_ram_0_0_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_ram_0_0_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_ram_0_0_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_ram_0_0_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_ram_0_1_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_ram_0_1_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_ram_0_1_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_ram_0_1_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_ram_0_2_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_ram_0_2_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_ram_0_2_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_ram_0_2_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_ram_0_3_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_ram_0_3_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_ram_0_3_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_ram_0_3_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_ram_0_4_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_ram_0_4_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_ram_0_4_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_ram_0_4_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_ram_0_5_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_ram_0_5_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_ram_0_5_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_ram_0_5_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_ram_0_6_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_ram_0_6_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_ram_0_6_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_ram_0_6_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  data_ram_0_7_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  data_ram_0_7_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  data_ram_0_7_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  data_ram_0_7_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  data_ram_1_0_0 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  data_ram_1_0_1 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  data_ram_1_0_2 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  data_ram_1_0_3 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  data_ram_1_1_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  data_ram_1_1_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  data_ram_1_1_2 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  data_ram_1_1_3 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  data_ram_1_2_0 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  data_ram_1_2_1 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  data_ram_1_2_2 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  data_ram_1_2_3 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  data_ram_1_3_0 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  data_ram_1_3_1 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  data_ram_1_3_2 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  data_ram_1_3_3 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  data_ram_1_4_0 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  data_ram_1_4_1 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  data_ram_1_4_2 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  data_ram_1_4_3 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  data_ram_1_5_0 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  data_ram_1_5_1 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  data_ram_1_5_2 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  data_ram_1_5_3 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  data_ram_1_6_0 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  data_ram_1_6_1 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  data_ram_1_6_2 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  data_ram_1_6_3 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  data_ram_1_7_0 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  data_ram_1_7_1 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  data_ram_1_7_2 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  data_ram_1_7_3 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  data_ram_2_0_0 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  data_ram_2_0_1 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  data_ram_2_0_2 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  data_ram_2_0_3 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  data_ram_2_1_0 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  data_ram_2_1_1 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  data_ram_2_1_2 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  data_ram_2_1_3 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  data_ram_2_2_0 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  data_ram_2_2_1 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  data_ram_2_2_2 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  data_ram_2_2_3 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  data_ram_2_3_0 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  data_ram_2_3_1 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  data_ram_2_3_2 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  data_ram_2_3_3 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  data_ram_2_4_0 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  data_ram_2_4_1 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  data_ram_2_4_2 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  data_ram_2_4_3 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  data_ram_2_5_0 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  data_ram_2_5_1 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  data_ram_2_5_2 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  data_ram_2_5_3 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  data_ram_2_6_0 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  data_ram_2_6_1 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  data_ram_2_6_2 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  data_ram_2_6_3 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  data_ram_2_7_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  data_ram_2_7_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  data_ram_2_7_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  data_ram_2_7_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  data_ram_3_0_0 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  data_ram_3_0_1 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  data_ram_3_0_2 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  data_ram_3_0_3 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  data_ram_3_1_0 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  data_ram_3_1_1 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  data_ram_3_1_2 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  data_ram_3_1_3 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  data_ram_3_2_0 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  data_ram_3_2_1 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  data_ram_3_2_2 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  data_ram_3_2_3 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  data_ram_3_3_0 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  data_ram_3_3_1 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  data_ram_3_3_2 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  data_ram_3_3_3 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  data_ram_3_4_0 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  data_ram_3_4_1 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  data_ram_3_4_2 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  data_ram_3_4_3 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  data_ram_3_5_0 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  data_ram_3_5_1 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  data_ram_3_5_2 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  data_ram_3_5_3 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  data_ram_3_6_0 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  data_ram_3_6_1 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  data_ram_3_6_2 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  data_ram_3_6_3 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  data_ram_3_7_0 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  data_ram_3_7_1 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  data_ram_3_7_2 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  data_ram_3_7_3 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  instrId_ram_0 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  instrId_ram_1 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  instrId_ram_2 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  instrId_ram_3 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  enqPtr = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  deqPtr = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  entryValid_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  entryValid_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  entryValid_2 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  entryValid_3 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  entryFrozen_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  entryFrozen_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  entryFrozen_2 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  entryFrozen_3 = _RAND_177[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_50(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_instrId,
  input  [31:0] io_enq_bits_data_0,
  input  [31:0] io_enq_bits_data_1,
  input  [31:0] io_enq_bits_data_2,
  input  [31:0] io_enq_bits_data_3,
  input  [31:0] io_enq_bits_data_4,
  input  [31:0] io_enq_bits_data_5,
  input  [31:0] io_enq_bits_data_6,
  input  [31:0] io_enq_bits_data_7,
  input         io_enq_bits_activeMask_0,
  input         io_enq_bits_activeMask_1,
  input         io_enq_bits_activeMask_2,
  input         io_enq_bits_activeMask_3,
  input         io_enq_bits_activeMask_4,
  input         io_enq_bits_activeMask_5,
  input         io_enq_bits_activeMask_6,
  input         io_enq_bits_activeMask_7,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_instrId,
  output [31:0] io_deq_bits_data_0,
  output [31:0] io_deq_bits_data_1,
  output [31:0] io_deq_bits_data_2,
  output [31:0] io_deq_bits_data_3,
  output [31:0] io_deq_bits_data_4,
  output [31:0] io_deq_bits_data_5,
  output [31:0] io_deq_bits_data_6,
  output [31:0] io_deq_bits_data_7,
  output        io_deq_bits_activeMask_0,
  output        io_deq_bits_activeMask_1,
  output        io_deq_bits_activeMask_2,
  output        io_deq_bits_activeMask_3,
  output        io_deq_bits_activeMask_4,
  output        io_deq_bits_activeMask_5,
  output        io_deq_bits_activeMask_6,
  output        io_deq_bits_activeMask_7,
  output [2:0]  io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_instrId [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_instrId_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_instrId_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_instrId_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_instrId_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_instrId_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_instrId_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_instrId_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_0 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_1 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_2 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_3 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_4 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_5 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_6 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_data_7 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_data_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_0 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_1 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_2 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_3 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_4 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_5 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_6 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_activeMask_7 [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_activeMask_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_activeMask_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire [1:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 312:32]
  wire [2:0] _io_count_T_1 = maybe_full & ptr_match ? 3'h4 : 3'h0; // @[Decoupled.scala 315:20]
  wire [2:0] _GEN_29 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 315:62]
  assign ram_instrId_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instrId_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instrId_io_deq_bits_MPORT_data = ram_instrId[ram_instrId_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_instrId_MPORT_data = io_enq_bits_instrId;
  assign ram_instrId_MPORT_addr = enq_ptr_value;
  assign ram_instrId_MPORT_mask = 1'h1;
  assign ram_instrId_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_0_io_deq_bits_MPORT_data = ram_data_0[ram_data_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_0_MPORT_data = io_enq_bits_data_0;
  assign ram_data_0_MPORT_addr = enq_ptr_value;
  assign ram_data_0_MPORT_mask = 1'h1;
  assign ram_data_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_1_io_deq_bits_MPORT_data = ram_data_1[ram_data_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_1_MPORT_data = io_enq_bits_data_1;
  assign ram_data_1_MPORT_addr = enq_ptr_value;
  assign ram_data_1_MPORT_mask = 1'h1;
  assign ram_data_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_2_io_deq_bits_MPORT_data = ram_data_2[ram_data_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_2_MPORT_data = io_enq_bits_data_2;
  assign ram_data_2_MPORT_addr = enq_ptr_value;
  assign ram_data_2_MPORT_mask = 1'h1;
  assign ram_data_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_3_io_deq_bits_MPORT_data = ram_data_3[ram_data_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_3_MPORT_data = io_enq_bits_data_3;
  assign ram_data_3_MPORT_addr = enq_ptr_value;
  assign ram_data_3_MPORT_mask = 1'h1;
  assign ram_data_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_4_io_deq_bits_MPORT_data = ram_data_4[ram_data_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_4_MPORT_data = io_enq_bits_data_4;
  assign ram_data_4_MPORT_addr = enq_ptr_value;
  assign ram_data_4_MPORT_mask = 1'h1;
  assign ram_data_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_5_io_deq_bits_MPORT_data = ram_data_5[ram_data_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_5_MPORT_data = io_enq_bits_data_5;
  assign ram_data_5_MPORT_addr = enq_ptr_value;
  assign ram_data_5_MPORT_mask = 1'h1;
  assign ram_data_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_6_io_deq_bits_MPORT_data = ram_data_6[ram_data_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_6_MPORT_data = io_enq_bits_data_6;
  assign ram_data_6_MPORT_addr = enq_ptr_value;
  assign ram_data_6_MPORT_mask = 1'h1;
  assign ram_data_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_7_io_deq_bits_MPORT_data = ram_data_7[ram_data_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_7_MPORT_data = io_enq_bits_data_7;
  assign ram_data_7_MPORT_addr = enq_ptr_value;
  assign ram_data_7_MPORT_mask = 1'h1;
  assign ram_data_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_0_io_deq_bits_MPORT_data = ram_activeMask_0[ram_activeMask_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_0_MPORT_data = io_enq_bits_activeMask_0;
  assign ram_activeMask_0_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_0_MPORT_mask = 1'h1;
  assign ram_activeMask_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_1_io_deq_bits_MPORT_data = ram_activeMask_1[ram_activeMask_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_1_MPORT_data = io_enq_bits_activeMask_1;
  assign ram_activeMask_1_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_1_MPORT_mask = 1'h1;
  assign ram_activeMask_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_2_io_deq_bits_MPORT_data = ram_activeMask_2[ram_activeMask_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_2_MPORT_data = io_enq_bits_activeMask_2;
  assign ram_activeMask_2_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_2_MPORT_mask = 1'h1;
  assign ram_activeMask_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_3_io_deq_bits_MPORT_data = ram_activeMask_3[ram_activeMask_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_3_MPORT_data = io_enq_bits_activeMask_3;
  assign ram_activeMask_3_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_3_MPORT_mask = 1'h1;
  assign ram_activeMask_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_4_io_deq_bits_MPORT_data = ram_activeMask_4[ram_activeMask_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_4_MPORT_data = io_enq_bits_activeMask_4;
  assign ram_activeMask_4_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_4_MPORT_mask = 1'h1;
  assign ram_activeMask_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_5_io_deq_bits_MPORT_data = ram_activeMask_5[ram_activeMask_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_5_MPORT_data = io_enq_bits_activeMask_5;
  assign ram_activeMask_5_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_5_MPORT_mask = 1'h1;
  assign ram_activeMask_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_6_io_deq_bits_MPORT_data = ram_activeMask_6[ram_activeMask_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_6_MPORT_data = io_enq_bits_activeMask_6;
  assign ram_activeMask_6_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_6_MPORT_mask = 1'h1;
  assign ram_activeMask_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_activeMask_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_activeMask_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_activeMask_7_io_deq_bits_MPORT_data = ram_activeMask_7[ram_activeMask_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_activeMask_7_MPORT_data = io_enq_bits_activeMask_7;
  assign ram_activeMask_7_MPORT_addr = enq_ptr_value;
  assign ram_activeMask_7_MPORT_mask = 1'h1;
  assign ram_activeMask_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_instrId = ram_instrId_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_0 = ram_data_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_1 = ram_data_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_2 = ram_data_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_3 = ram_data_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_4 = ram_data_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_5 = ram_data_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_6 = ram_data_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data_7 = ram_data_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_0 = ram_activeMask_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_1 = ram_activeMask_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_2 = ram_activeMask_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_3 = ram_activeMask_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_4 = ram_activeMask_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_5 = ram_activeMask_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_6 = ram_activeMask_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_activeMask_7 = ram_activeMask_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_count = _io_count_T_1 | _GEN_29; // @[Decoupled.scala 315:62]
  always @(posedge clock) begin
    if (ram_instrId_MPORT_en & ram_instrId_MPORT_mask) begin
      ram_instrId[ram_instrId_MPORT_addr] <= ram_instrId_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_0_MPORT_en & ram_data_0_MPORT_mask) begin
      ram_data_0[ram_data_0_MPORT_addr] <= ram_data_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_1_MPORT_en & ram_data_1_MPORT_mask) begin
      ram_data_1[ram_data_1_MPORT_addr] <= ram_data_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_2_MPORT_en & ram_data_2_MPORT_mask) begin
      ram_data_2[ram_data_2_MPORT_addr] <= ram_data_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_3_MPORT_en & ram_data_3_MPORT_mask) begin
      ram_data_3[ram_data_3_MPORT_addr] <= ram_data_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_4_MPORT_en & ram_data_4_MPORT_mask) begin
      ram_data_4[ram_data_4_MPORT_addr] <= ram_data_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_5_MPORT_en & ram_data_5_MPORT_mask) begin
      ram_data_5[ram_data_5_MPORT_addr] <= ram_data_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_6_MPORT_en & ram_data_6_MPORT_mask) begin
      ram_data_6[ram_data_6_MPORT_addr] <= ram_data_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_7_MPORT_en & ram_data_7_MPORT_mask) begin
      ram_data_7[ram_data_7_MPORT_addr] <= ram_data_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_0_MPORT_en & ram_activeMask_0_MPORT_mask) begin
      ram_activeMask_0[ram_activeMask_0_MPORT_addr] <= ram_activeMask_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_1_MPORT_en & ram_activeMask_1_MPORT_mask) begin
      ram_activeMask_1[ram_activeMask_1_MPORT_addr] <= ram_activeMask_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_2_MPORT_en & ram_activeMask_2_MPORT_mask) begin
      ram_activeMask_2[ram_activeMask_2_MPORT_addr] <= ram_activeMask_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_3_MPORT_en & ram_activeMask_3_MPORT_mask) begin
      ram_activeMask_3[ram_activeMask_3_MPORT_addr] <= ram_activeMask_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_4_MPORT_en & ram_activeMask_4_MPORT_mask) begin
      ram_activeMask_4[ram_activeMask_4_MPORT_addr] <= ram_activeMask_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_5_MPORT_en & ram_activeMask_5_MPORT_mask) begin
      ram_activeMask_5[ram_activeMask_5_MPORT_addr] <= ram_activeMask_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_6_MPORT_en & ram_activeMask_6_MPORT_mask) begin
      ram_activeMask_6[ram_activeMask_6_MPORT_addr] <= ram_activeMask_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_activeMask_7_MPORT_en & ram_activeMask_7_MPORT_mask) begin
      ram_activeMask_7[ram_activeMask_7_MPORT_addr] <= ram_activeMask_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instrId[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_0[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_1[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_2[initvar] = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_3[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_4[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_5[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_6[initvar] = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data_7[initvar] = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_0[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_1[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_2[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_3[initvar] = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_4[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_5[initvar] = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_6[initvar] = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_activeMask_7[initvar] = _RAND_16[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  enq_ptr_value = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  deq_ptr_value = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  maybe_full = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_3(
  input        clock,
  input        reset,
  input        io_r_req_valid,
  input  [5:0] io_r_req_bits_setIdx,
  output [7:0] io_r_resp_data_0,
  output [7:0] io_r_resp_data_1,
  output [7:0] io_r_resp_data_2,
  output [7:0] io_r_resp_data_3,
  input        io_w_req_valid,
  input  [5:0] io_w_req_bits_setIdx,
  input  [7:0] io_w_req_bits_data_0,
  input  [7:0] io_w_req_bits_data_1,
  input  [7:0] io_w_req_bits_data_2,
  input  [7:0] io_w_req_bits_data_3,
  input  [3:0] io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] array_0 [0:63]; // @[SRAMTemplate.scala 101:26]
  wire  array_0_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_0_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_0_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_0_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_0_raw_rdata_en_pipe_0;
  reg [5:0] array_0_raw_rdata_addr_pipe_0;
  reg [7:0] array_1 [0:63]; // @[SRAMTemplate.scala 101:26]
  wire  array_1_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_1_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_1_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_1_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_1_raw_rdata_en_pipe_0;
  reg [5:0] array_1_raw_rdata_addr_pipe_0;
  reg [7:0] array_2 [0:63]; // @[SRAMTemplate.scala 101:26]
  wire  array_2_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_2_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_2_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_2_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_2_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_2_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_2_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_2_raw_rdata_en_pipe_0;
  reg [5:0] array_2_raw_rdata_addr_pipe_0;
  reg [7:0] array_3 [0:63]; // @[SRAMTemplate.scala 101:26]
  wire  array_3_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_3_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_3_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_3_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [5:0] array_3_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_3_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_3_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_3_raw_rdata_en_pipe_0;
  reg [5:0] array_3_raw_rdata_addr_pipe_0;
  reg [63:0] bypass_wdata_lfsr; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor = bypass_wdata_lfsr[0] ^ bypass_wdata_lfsr[1] ^ bypass_wdata_lfsr[3] ^ bypass_wdata_lfsr[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_2 = {bypass_wdata_xor,bypass_wdata_lfsr[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_1; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_1 = bypass_wdata_lfsr_1[0] ^ bypass_wdata_lfsr_1[1] ^ bypass_wdata_lfsr_1[3] ^
    bypass_wdata_lfsr_1[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_6 = {bypass_wdata_xor_1,bypass_wdata_lfsr_1[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_2; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_2 = bypass_wdata_lfsr_2[0] ^ bypass_wdata_lfsr_2[1] ^ bypass_wdata_lfsr_2[3] ^
    bypass_wdata_lfsr_2[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_10 = {bypass_wdata_xor_2,bypass_wdata_lfsr_2[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_3; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_3 = bypass_wdata_lfsr_3[0] ^ bypass_wdata_lfsr_3[1] ^ bypass_wdata_lfsr_3[3] ^
    bypass_wdata_lfsr_3[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_14 = {bypass_wdata_xor_3,bypass_wdata_lfsr_3[63:1]}; // @[Cat.scala 31:58]
  reg  bypass_mask_need_check; // @[SRAMTemplate.scala 126:29]
  reg [5:0] bypass_mask_waddr_reg; // @[SRAMTemplate.scala 127:28]
  reg [5:0] bypass_mask_raddr_reg; // @[SRAMTemplate.scala 128:28]
  wire  _bypass_mask_bypass_T_1 = bypass_mask_need_check & bypass_mask_waddr_reg == bypass_mask_raddr_reg; // @[SRAMTemplate.scala 130:39]
  wire [3:0] _bypass_mask_bypass_T_3 = _bypass_mask_bypass_T_1 ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  reg [3:0] bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:76]
  wire [3:0] bypass_mask_bypass = _bypass_mask_bypass_T_3 & bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:67]
  wire [7:0] bypass_wdata_0 = bypass_wdata_lfsr[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [7:0] bypass_wdata_1 = bypass_wdata_lfsr_1[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [7:0] bypass_wdata_2 = bypass_wdata_lfsr_2[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [7:0] bypass_wdata_3 = bypass_wdata_lfsr_3[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  assign array_0_raw_rdata_en = array_0_raw_rdata_en_pipe_0;
  assign array_0_raw_rdata_addr = array_0_raw_rdata_addr_pipe_0;
  assign array_0_raw_rdata_data = array_0[array_0_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_0_MPORT_data = io_w_req_bits_data_0;
  assign array_0_MPORT_addr = io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = io_w_req_bits_waymask[0];
  assign array_0_MPORT_en = io_w_req_valid;
  assign array_1_raw_rdata_en = array_1_raw_rdata_en_pipe_0;
  assign array_1_raw_rdata_addr = array_1_raw_rdata_addr_pipe_0;
  assign array_1_raw_rdata_data = array_1[array_1_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_1_MPORT_data = io_w_req_bits_data_1;
  assign array_1_MPORT_addr = io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = io_w_req_bits_waymask[1];
  assign array_1_MPORT_en = io_w_req_valid;
  assign array_2_raw_rdata_en = array_2_raw_rdata_en_pipe_0;
  assign array_2_raw_rdata_addr = array_2_raw_rdata_addr_pipe_0;
  assign array_2_raw_rdata_data = array_2[array_2_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_2_MPORT_data = io_w_req_bits_data_2;
  assign array_2_MPORT_addr = io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = io_w_req_bits_waymask[2];
  assign array_2_MPORT_en = io_w_req_valid;
  assign array_3_raw_rdata_en = array_3_raw_rdata_en_pipe_0;
  assign array_3_raw_rdata_addr = array_3_raw_rdata_addr_pipe_0;
  assign array_3_raw_rdata_data = array_3[array_3_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_3_MPORT_data = io_w_req_bits_data_3;
  assign array_3_MPORT_addr = io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = io_w_req_bits_waymask[3];
  assign array_3_MPORT_en = io_w_req_valid;
  assign io_r_resp_data_0 = bypass_mask_bypass[0] ? bypass_wdata_0 : array_0_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_1 = bypass_mask_bypass[1] ? bypass_wdata_1 : array_1_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_2 = bypass_mask_bypass[2] ? bypass_wdata_2 : array_2_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_3 = bypass_mask_bypass[3] ? bypass_wdata_3 : array_3_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_0_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_0_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_1_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_1_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_2_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_2_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_3_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_3_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr <= 64'h1;
    end else begin
      bypass_wdata_lfsr <= _bypass_wdata_lfsr_T_2;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_1 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_1 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_1 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_1 <= _bypass_wdata_lfsr_T_6;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_2 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_2 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_2 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_2 <= _bypass_wdata_lfsr_T_10;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_3 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_3 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_3 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_3 <= _bypass_wdata_lfsr_T_14;
    end
    bypass_mask_need_check <= io_r_req_valid & io_w_req_valid; // @[SRAMTemplate.scala 126:34]
    bypass_mask_waddr_reg <= io_w_req_bits_setIdx; // @[SRAMTemplate.scala 127:28]
    bypass_mask_raddr_reg <= io_r_req_bits_setIdx; // @[SRAMTemplate.scala 128:28]
    bypass_mask_bypass_REG <= io_w_req_bits_waymask; // @[SRAMTemplate.scala 130:76]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    array_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    array_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    array_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    array_3[initvar] = _RAND_9[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_raw_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_raw_rdata_addr_pipe_0 = _RAND_2[5:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_raw_rdata_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_raw_rdata_addr_pipe_0 = _RAND_5[5:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_raw_rdata_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_raw_rdata_addr_pipe_0 = _RAND_8[5:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_raw_rdata_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_raw_rdata_addr_pipe_0 = _RAND_11[5:0];
  _RAND_12 = {2{`RANDOM}};
  bypass_wdata_lfsr = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  bypass_wdata_lfsr_1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  bypass_wdata_lfsr_2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  bypass_wdata_lfsr_3 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  bypass_mask_need_check = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  bypass_mask_waddr_reg = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  bypass_mask_raddr_reg = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  bypass_mask_bypass_REG = _RAND_19[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_15(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_a_source,
  input  [31:0] io_in_0_bits_a_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [2:0]  io_in_1_bits_a_opcode,
  input  [1:0]  io_in_1_bits_a_source,
  input  [31:0] io_in_1_bits_a_addr,
  input  [31:0] io_in_1_bits_a_data_0,
  input  [31:0] io_in_1_bits_a_data_1,
  input  [31:0] io_in_1_bits_a_data_2,
  input  [31:0] io_in_1_bits_a_data_3,
  input  [31:0] io_in_1_bits_a_data_4,
  input  [31:0] io_in_1_bits_a_data_5,
  input  [31:0] io_in_1_bits_a_data_6,
  input  [31:0] io_in_1_bits_a_data_7,
  input         io_in_1_bits_a_mask_0,
  input         io_in_1_bits_a_mask_1,
  input         io_in_1_bits_a_mask_2,
  input         io_in_1_bits_a_mask_3,
  input         io_in_1_bits_a_mask_4,
  input         io_in_1_bits_a_mask_5,
  input         io_in_1_bits_a_mask_6,
  input         io_in_1_bits_a_mask_7,
  input         io_out_ready,
  output        io_out_valid,
  output [2:0]  io_out_bits_a_opcode,
  output [1:0]  io_out_bits_a_source,
  output [31:0] io_out_bits_a_addr,
  output [31:0] io_out_bits_a_data_0,
  output [31:0] io_out_bits_a_data_1,
  output [31:0] io_out_bits_a_data_2,
  output [31:0] io_out_bits_a_data_3,
  output [31:0] io_out_bits_a_data_4,
  output [31:0] io_out_bits_a_data_5,
  output [31:0] io_out_bits_a_data_6,
  output [31:0] io_out_bits_a_data_7,
  output        io_out_bits_a_mask_0,
  output        io_out_bits_a_mask_1,
  output        io_out_bits_a_mask_2,
  output        io_out_bits_a_mask_3,
  output        io_out_bits_a_mask_4,
  output        io_out_bits_a_mask_5,
  output        io_out_bits_a_mask_6,
  output        io_out_bits_a_mask_7
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_a_opcode = io_in_0_valid ? 3'h4 : io_in_1_bits_a_opcode; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_source = io_in_0_valid ? io_in_0_bits_a_source : io_in_1_bits_a_source; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_addr = io_in_0_valid ? io_in_0_bits_a_addr : io_in_1_bits_a_addr; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_0 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_0; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_1 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_1; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_2 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_2; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_3 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_3; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_4 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_4; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_5 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_5; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_6 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_6; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_data_7 = io_in_0_valid ? 32'h0 : io_in_1_bits_a_data_7; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_0 = io_in_0_valid | io_in_1_bits_a_mask_0; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_1 = io_in_0_valid | io_in_1_bits_a_mask_1; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_2 = io_in_0_valid | io_in_1_bits_a_mask_2; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_3 = io_in_0_valid | io_in_1_bits_a_mask_3; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_4 = io_in_0_valid | io_in_1_bits_a_mask_4; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_5 = io_in_0_valid | io_in_1_bits_a_mask_5; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_6 = io_in_0_valid | io_in_1_bits_a_mask_6; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_a_mask_7 = io_in_0_valid | io_in_1_bits_a_mask_7; // @[Arbiter.scala 139:15 141:26 143:19]
endmodule
module DataCache(
  input         clock,
  input         reset,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [1:0]  io_coreReq_bits_instrId,
  input         io_coreReq_bits_isWrite,
  input  [21:0] io_coreReq_bits_tag,
  input  [4:0]  io_coreReq_bits_setIdx,
  input         io_coreReq_bits_perLaneAddr_0_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_0_blockOffset,
  input         io_coreReq_bits_perLaneAddr_1_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_1_blockOffset,
  input         io_coreReq_bits_perLaneAddr_2_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_2_blockOffset,
  input         io_coreReq_bits_perLaneAddr_3_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_3_blockOffset,
  input         io_coreReq_bits_perLaneAddr_4_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_4_blockOffset,
  input         io_coreReq_bits_perLaneAddr_5_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_5_blockOffset,
  input         io_coreReq_bits_perLaneAddr_6_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_6_blockOffset,
  input         io_coreReq_bits_perLaneAddr_7_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_7_blockOffset,
  input  [31:0] io_coreReq_bits_data_0,
  input  [31:0] io_coreReq_bits_data_1,
  input  [31:0] io_coreReq_bits_data_2,
  input  [31:0] io_coreReq_bits_data_3,
  input  [31:0] io_coreReq_bits_data_4,
  input  [31:0] io_coreReq_bits_data_5,
  input  [31:0] io_coreReq_bits_data_6,
  input  [31:0] io_coreReq_bits_data_7,
  input         io_coreRsp_ready,
  output        io_coreRsp_valid,
  output [1:0]  io_coreRsp_bits_instrId,
  output [31:0] io_coreRsp_bits_data_0,
  output [31:0] io_coreRsp_bits_data_1,
  output [31:0] io_coreRsp_bits_data_2,
  output [31:0] io_coreRsp_bits_data_3,
  output [31:0] io_coreRsp_bits_data_4,
  output [31:0] io_coreRsp_bits_data_5,
  output [31:0] io_coreRsp_bits_data_6,
  output [31:0] io_coreRsp_bits_data_7,
  output        io_coreRsp_bits_activeMask_0,
  output        io_coreRsp_bits_activeMask_1,
  output        io_coreRsp_bits_activeMask_2,
  output        io_coreRsp_bits_activeMask_3,
  output        io_coreRsp_bits_activeMask_4,
  output        io_coreRsp_bits_activeMask_5,
  output        io_coreRsp_bits_activeMask_6,
  output        io_coreRsp_bits_activeMask_7,
  output        io_memRsp_ready,
  input         io_memRsp_valid,
  input  [31:0] io_memRsp_bits_d_addr,
  input  [31:0] io_memRsp_bits_d_data_0,
  input  [31:0] io_memRsp_bits_d_data_1,
  input  [31:0] io_memRsp_bits_d_data_2,
  input  [31:0] io_memRsp_bits_d_data_3,
  input  [31:0] io_memRsp_bits_d_data_4,
  input  [31:0] io_memRsp_bits_d_data_5,
  input  [31:0] io_memRsp_bits_d_data_6,
  input  [31:0] io_memRsp_bits_d_data_7,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [2:0]  io_memReq_bits_a_opcode,
  output [1:0]  io_memReq_bits_a_source,
  output [31:0] io_memReq_bits_a_addr,
  output [31:0] io_memReq_bits_a_data_0,
  output [31:0] io_memReq_bits_a_data_1,
  output [31:0] io_memReq_bits_a_data_2,
  output [31:0] io_memReq_bits_a_data_3,
  output [31:0] io_memReq_bits_a_data_4,
  output [31:0] io_memReq_bits_a_data_5,
  output [31:0] io_memReq_bits_a_data_6,
  output [31:0] io_memReq_bits_a_data_7,
  output        io_memReq_bits_a_mask_0,
  output        io_memReq_bits_a_mask_1,
  output        io_memReq_bits_a_mask_2,
  output        io_memReq_bits_a_mask_3,
  output        io_memReq_bits_a_mask_4,
  output        io_memReq_bits_a_mask_5,
  output        io_memReq_bits_a_mask_6,
  output        io_memReq_bits_a_mask_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
`endif // RANDOMIZE_REG_INIT
  wire  BankConfArb_clock; // @[DCache.scala 85:27]
  wire  BankConfArb_reset; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_isWrite; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_enable; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_0_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_0_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_0_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_1_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_1_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_1_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_2_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_2_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_2_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_3_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_3_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_3_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_4_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_4_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_4_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_5_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_5_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_5_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_6_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_6_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_6_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_7_activeMask; // @[DCache.scala 85:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_7_blockOffset; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_coreReqArb_perLaneAddr_7_wordOffset1H; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_0; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_1; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_2; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_3; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_4; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_5; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_6; // @[DCache.scala 85:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_7; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_0_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_1_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_2_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_3_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_4_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_5_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_6_wordOffset1H; // @[DCache.scala 85:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_7_wordOffset1H; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_0; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_1; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_2; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_3; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_4; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_5; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_6; // @[DCache.scala 85:27]
  wire  BankConfArb_io_dataArrayEn_7; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_0; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_1; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_2; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_3; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_4; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_5; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_6; // @[DCache.scala 85:27]
  wire  BankConfArb_io_activeLane_7; // @[DCache.scala 85:27]
  wire  BankConfArb_io_bankConflict; // @[DCache.scala 85:27]
  wire  MshrAccess_clock; // @[DCache.scala 87:26]
  wire  MshrAccess_reset; // @[DCache.scala 87:26]
  wire  MshrAccess_io_missReq_ready; // @[DCache.scala 87:26]
  wire  MshrAccess_io_missReq_valid; // @[DCache.scala 87:26]
  wire [26:0] MshrAccess_io_missReq_bits_blockAddr; // @[DCache.scala 87:26]
  wire [1:0] MshrAccess_io_missReq_bits_instrId; // @[DCache.scala 87:26]
  wire [64:0] MshrAccess_io_missReq_bits_targetInfo; // @[DCache.scala 87:26]
  wire  MshrAccess_io_missRspIn_ready; // @[DCache.scala 87:26]
  wire  MshrAccess_io_missRspIn_valid; // @[DCache.scala 87:26]
  wire [26:0] MshrAccess_io_missRspIn_bits_blockAddr; // @[DCache.scala 87:26]
  wire  MshrAccess_io_missRspOut_ready; // @[DCache.scala 87:26]
  wire  MshrAccess_io_missRspOut_valid; // @[DCache.scala 87:26]
  wire [64:0] MshrAccess_io_missRspOut_bits_targetInfo; // @[DCache.scala 87:26]
  wire [26:0] MshrAccess_io_missRspOut_bits_blockAddr; // @[DCache.scala 87:26]
  wire [1:0] MshrAccess_io_missRspOut_bits_instrId; // @[DCache.scala 87:26]
  wire  MshrAccess_io_miss2mem_ready; // @[DCache.scala 87:26]
  wire  MshrAccess_io_miss2mem_valid; // @[DCache.scala 87:26]
  wire [26:0] MshrAccess_io_miss2mem_bits_blockAddr; // @[DCache.scala 87:26]
  wire [1:0] MshrAccess_io_miss2mem_bits_instrId; // @[DCache.scala 87:26]
  wire  TagAccess_clock; // @[DCache.scala 90:25]
  wire  TagAccess_reset; // @[DCache.scala 90:25]
  wire  TagAccess_io_r_req_valid; // @[DCache.scala 90:25]
  wire [4:0] TagAccess_io_r_req_bits_setIdx; // @[DCache.scala 90:25]
  wire [21:0] TagAccess_io_tagFromCore_st1; // @[DCache.scala 90:25]
  wire  TagAccess_io_coreReqReady; // @[DCache.scala 90:25]
  wire  TagAccess_io_w_req_valid; // @[DCache.scala 90:25]
  wire [4:0] TagAccess_io_w_req_bits_setIdx; // @[DCache.scala 90:25]
  wire [21:0] TagAccess_io_w_req_bits_data_0; // @[DCache.scala 90:25]
  wire [21:0] TagAccess_io_w_req_bits_data_1; // @[DCache.scala 90:25]
  wire [1:0] TagAccess_io_waymaskReplacement; // @[DCache.scala 90:25]
  wire [1:0] TagAccess_io_waymaskHit_st1; // @[DCache.scala 90:25]
  wire  TagAccess_io_hit_st1; // @[DCache.scala 90:25]
  wire [31:0] DataCorssBar_io_DataIn_0; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_1; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_2; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_3; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_4; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_5; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_6; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataIn_7; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_0; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_1; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_2; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_3; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_4; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_5; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_6; // @[DCache.scala 91:28]
  wire [31:0] DataCorssBar_io_DataOut_7; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_0; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_1; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_2; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_3; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_4; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_5; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_6; // @[DCache.scala 91:28]
  wire [7:0] DataCorssBar_io_Select1H_7; // @[DCache.scala 91:28]
  wire  WriteDataBuf_clock; // @[DCache.scala 92:28]
  wire  WriteDataBuf_reset; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_inputBus_ready; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_inputBus_valid; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_0; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_1; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_2; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_3; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_4; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_5; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_6; // @[DCache.scala 92:28]
  wire [3:0] WriteDataBuf_io_inputBus_bits_mask_7; // @[DCache.scala 92:28]
  wire [31:0] WriteDataBuf_io_inputBus_bits_addr; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_0_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_0_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_0_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_0_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_1_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_1_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_1_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_1_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_2_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_2_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_2_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_2_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_3_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_3_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_3_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_3_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_4_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_4_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_4_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_4_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_5_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_5_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_5_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_5_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_6_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_6_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_6_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_6_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_7_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_7_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_7_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_inputBus_bits_data_7_3; // @[DCache.scala 92:28]
  wire [1:0] WriteDataBuf_io_inputBus_bits_instrId; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_inputBus_bits_bankConflict; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_inputBus_bits_subWordMissReq; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_inputBus_bits_subWordMissRsp; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_ready; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_valid; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_0; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_1; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_2; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_3; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_4; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_5; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_6; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_outputBus_bits_mask_7; // @[DCache.scala 92:28]
  wire [31:0] WriteDataBuf_io_outputBus_bits_addr; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_0_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_0_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_0_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_0_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_1_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_1_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_1_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_1_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_2_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_2_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_2_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_2_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_3_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_3_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_3_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_3_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_4_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_4_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_4_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_4_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_5_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_5_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_5_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_5_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_6_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_6_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_6_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_6_3; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_7_0; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_7_1; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_7_2; // @[DCache.scala 92:28]
  wire [7:0] WriteDataBuf_io_outputBus_bits_data_7_3; // @[DCache.scala 92:28]
  wire [1:0] WriteDataBuf_io_outputBus_bits_instrId; // @[DCache.scala 92:28]
  wire  WriteDataBuf_io_wdbAlmostFull; // @[DCache.scala 92:28]
  wire  coreRsp_Q_clock; // @[DCache.scala 96:25]
  wire  coreRsp_Q_reset; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_ready; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_valid; // @[DCache.scala 96:25]
  wire [1:0] coreRsp_Q_io_enq_bits_instrId; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_0; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_1; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_2; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_3; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_4; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_5; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_6; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_7; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_0; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_1; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_2; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_3; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_4; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_5; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_6; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_7; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_ready; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_valid; // @[DCache.scala 96:25]
  wire [1:0] coreRsp_Q_io_deq_bits_instrId; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_0; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_1; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_2; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_3; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_4; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_5; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_6; // @[DCache.scala 96:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_7; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_0; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_1; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_2; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_3; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_4; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_5; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_6; // @[DCache.scala 96:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_7; // @[DCache.scala 96:25]
  wire [2:0] coreRsp_Q_io_count; // @[DCache.scala 96:25]
  wire  memRsp_Q_clock; // @[DCache.scala 99:24]
  wire  memRsp_Q_reset; // @[DCache.scala 99:24]
  wire  memRsp_Q_io_enq_ready; // @[DCache.scala 99:24]
  wire  memRsp_Q_io_enq_valid; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_addr; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_0; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_1; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_2; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_3; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_4; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_5; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_6; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_enq_bits_d_data_7; // @[DCache.scala 99:24]
  wire  memRsp_Q_io_deq_ready; // @[DCache.scala 99:24]
  wire  memRsp_Q_io_deq_valid; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_addr; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_0; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_1; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_2; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_3; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_4; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_5; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_6; // @[DCache.scala 99:24]
  wire [31:0] memRsp_Q_io_deq_bits_d_data_7; // @[DCache.scala 99:24]
  wire  DataAccessesRRsp_DataAccess_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_1_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_1_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_1_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_1_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_1_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_2_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_2_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_2_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_2_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_2_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_3_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_3_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_3_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_3_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_3_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_4_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_4_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_4_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_4_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_4_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_5_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_5_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_5_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_5_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_5_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_6_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_6_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_6_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_6_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_6_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_7_clock; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_7_reset; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_7_io_r_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_7_io_r_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_3; // @[DCache.scala 240:28]
  wire  DataAccessesRRsp_DataAccess_7_io_w_req_valid; // @[DCache.scala 240:28]
  wire [5:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_setIdx; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_0; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_1; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_2; // @[DCache.scala 240:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_3; // @[DCache.scala 240:28]
  wire [3:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_waymask; // @[DCache.scala 240:28]
  wire  MemReqArb_io_in_0_ready; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_0_valid; // @[DCache.scala 381:25]
  wire [1:0] MemReqArb_io_in_0_bits_a_source; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_0_bits_a_addr; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_ready; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_valid; // @[DCache.scala 381:25]
  wire [2:0] MemReqArb_io_in_1_bits_a_opcode; // @[DCache.scala 381:25]
  wire [1:0] MemReqArb_io_in_1_bits_a_source; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_addr; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_0; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_1; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_2; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_3; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_4; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_5; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_6; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_in_1_bits_a_data_7; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_0; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_1; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_2; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_3; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_4; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_5; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_6; // @[DCache.scala 381:25]
  wire  MemReqArb_io_in_1_bits_a_mask_7; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_ready; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_valid; // @[DCache.scala 381:25]
  wire [2:0] MemReqArb_io_out_bits_a_opcode; // @[DCache.scala 381:25]
  wire [1:0] MemReqArb_io_out_bits_a_source; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_addr; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_0; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_1; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_2; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_3; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_4; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_5; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_6; // @[DCache.scala 381:25]
  wire [31:0] MemReqArb_io_out_bits_a_data_7; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_0; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_1; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_2; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_3; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_4; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_5; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_6; // @[DCache.scala 381:25]
  wire  MemReqArb_io_out_bits_a_mask_7; // @[DCache.scala 381:25]
  wire  _coreReq_st1_T = io_coreReq_ready & io_coreReq_valid; // @[Decoupled.scala 50:35]
  reg [1:0] coreReq_st1_instrId; // @[Reg.scala 16:16]
  reg  coreReq_st1_isWrite; // @[Reg.scala 16:16]
  reg [21:0] coreReq_st1_tag; // @[Reg.scala 16:16]
  reg [4:0] coreReq_st1_setIdx; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_0_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_0_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_1_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_1_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_2_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_2_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_3_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_3_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_4_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_4_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_5_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_5_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_6_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_6_blockOffset; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_7_activeMask; // @[Reg.scala 16:16]
  reg [2:0] coreReq_st1_perLaneAddr_7_blockOffset; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_0; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_1; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_2; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_3; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_4; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_5; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_6; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_7; // @[Reg.scala 16:16]
  reg [1:0] coreReq_st2_instrId; // @[DCache.scala 105:28]
  reg  coreReq_st2_isWrite; // @[DCache.scala 105:28]
  reg [21:0] coreReq_st2_tag; // @[DCache.scala 105:28]
  reg [4:0] coreReq_st2_setIdx; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_0; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_1; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_2; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_3; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_4; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_5; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_6; // @[DCache.scala 105:28]
  reg [31:0] coreReq_st2_data_7; // @[DCache.scala 105:28]
  reg [1:0] coreReqInstrId_st3; // @[DCache.scala 106:35]
  reg  coreReqActvMask_st3_r_0; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_1; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_2; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_3; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_4; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_5; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_6; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_r_7; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_0; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_1; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_2; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_3; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_4; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_5; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_6; // @[Reg.scala 16:16]
  reg  coreReqActvMask_st3_7; // @[Reg.scala 16:16]
  wire  missRspFromMshr_st1 = MshrAccess_io_missRspOut_valid; // @[DCache.scala 204:23 88:33]
  wire [64:0] _missRspTI_st1_WIRE_1 = MshrAccess_io_missRspOut_bits_targetInfo;
  wire  missRspTI_st1_isWrite = _missRspTI_st1_WIRE_1[64]; // @[DCache.scala 205:69]
  reg  cacheHit_st1_REG; // @[DCache.scala 140:50]
  wire  cacheHit_st1 = TagAccess_io_hit_st1 & cacheHit_st1_REG; // @[DCache.scala 140:40]
  wire  missRspTI_st1_perLaneAddr_0_activeMask = _missRspTI_st1_WIRE_1[7]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_0_blockOffset = _missRspTI_st1_WIRE_1[6:4]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_0_wordOffset1H = _missRspTI_st1_WIRE_1[3:0]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_1_activeMask = _missRspTI_st1_WIRE_1[15]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_1_blockOffset = _missRspTI_st1_WIRE_1[14:12]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_1_wordOffset1H = _missRspTI_st1_WIRE_1[11:8]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_2_activeMask = _missRspTI_st1_WIRE_1[23]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_2_blockOffset = _missRspTI_st1_WIRE_1[22:20]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_2_wordOffset1H = _missRspTI_st1_WIRE_1[19:16]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_3_activeMask = _missRspTI_st1_WIRE_1[31]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_3_blockOffset = _missRspTI_st1_WIRE_1[30:28]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_3_wordOffset1H = _missRspTI_st1_WIRE_1[27:24]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_4_activeMask = _missRspTI_st1_WIRE_1[39]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_4_blockOffset = _missRspTI_st1_WIRE_1[38:36]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_4_wordOffset1H = _missRspTI_st1_WIRE_1[35:32]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_5_activeMask = _missRspTI_st1_WIRE_1[47]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_5_blockOffset = _missRspTI_st1_WIRE_1[46:44]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_5_wordOffset1H = _missRspTI_st1_WIRE_1[43:40]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_6_activeMask = _missRspTI_st1_WIRE_1[55]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_6_blockOffset = _missRspTI_st1_WIRE_1[54:52]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_6_wordOffset1H = _missRspTI_st1_WIRE_1[51:48]; // @[DCache.scala 205:69]
  wire  missRspTI_st1_perLaneAddr_7_activeMask = _missRspTI_st1_WIRE_1[63]; // @[DCache.scala 205:69]
  wire [2:0] missRspTI_st1_perLaneAddr_7_blockOffset = _missRspTI_st1_WIRE_1[62:60]; // @[DCache.scala 205:69]
  wire [3:0] missRspTI_st1_perLaneAddr_7_wordOffset1H = _missRspTI_st1_WIRE_1[59:56]; // @[DCache.scala 205:69]
  reg  cacheMiss_st1_r; // @[Reg.scala 16:16]
  wire  cacheMiss_st1 = ~TagAccess_io_hit_st1 & cacheMiss_st1_r; // @[DCache.scala 141:45]
  wire  wayIdxAtHit_st1 = TagAccess_io_waymaskHit_st1[1]; // @[CircuitMath.scala 30:8]
  reg  wayIdxAtHit_st2; // @[DCache.scala 145:32]
  wire  wayIdxReplace_st0 = TagAccess_io_waymaskReplacement[1]; // @[CircuitMath.scala 30:8]
  wire  _writeFullWordBank_st1_T = &BankConfArb_io_addrCrsbarOut_0_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_1 = &BankConfArb_io_addrCrsbarOut_1_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_2 = &BankConfArb_io_addrCrsbarOut_2_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_3 = &BankConfArb_io_addrCrsbarOut_3_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_4 = &BankConfArb_io_addrCrsbarOut_4_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_5 = &BankConfArb_io_addrCrsbarOut_5_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_6 = &BankConfArb_io_addrCrsbarOut_6_wordOffset1H; // @[DCache.scala 149:83]
  wire  _writeFullWordBank_st1_T_7 = &BankConfArb_io_addrCrsbarOut_7_wordOffset1H; // @[DCache.scala 149:83]
  wire [7:0] writeFullWordBank_st1 = {_writeFullWordBank_st1_T,_writeFullWordBank_st1_T_1,_writeFullWordBank_st1_T_2,
    _writeFullWordBank_st1_T_3,_writeFullWordBank_st1_T_4,_writeFullWordBank_st1_T_5,_writeFullWordBank_st1_T_6,
    _writeFullWordBank_st1_T_7}; // @[Cat.scala 31:58]
  wire  _writeTouchBank_st1_T = |BankConfArb_io_addrCrsbarOut_0_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_1 = |BankConfArb_io_addrCrsbarOut_1_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_2 = |BankConfArb_io_addrCrsbarOut_2_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_3 = |BankConfArb_io_addrCrsbarOut_3_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_4 = |BankConfArb_io_addrCrsbarOut_4_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_5 = |BankConfArb_io_addrCrsbarOut_5_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_6 = |BankConfArb_io_addrCrsbarOut_6_wordOffset1H; // @[DCache.scala 150:83]
  wire  _writeTouchBank_st1_T_7 = |BankConfArb_io_addrCrsbarOut_7_wordOffset1H; // @[DCache.scala 150:83]
  wire [7:0] writeTouchBank_st1 = {_writeTouchBank_st1_T,_writeTouchBank_st1_T_1,_writeTouchBank_st1_T_2,
    _writeTouchBank_st1_T_3,_writeTouchBank_st1_T_4,_writeTouchBank_st1_T_5,_writeTouchBank_st1_T_6,
    _writeTouchBank_st1_T_7}; // @[Cat.scala 31:58]
  wire [7:0] writeSubWordBank_st1 = writeFullWordBank_st1 ^ writeTouchBank_st1; // @[DCache.scala 151:52]
  wire  byteEn_st1 = writeFullWordBank_st1 != writeTouchBank_st1; // @[DCache.scala 152:49]
  wire  _readHit_st1_T = ~coreReq_st1_isWrite; // @[DCache.scala 154:36]
  wire  readHit_st1 = cacheHit_st1 & ~coreReq_st1_isWrite; // @[DCache.scala 154:34]
  wire  writeHit_st1 = cacheHit_st1 & coreReq_st1_isWrite; // @[DCache.scala 155:35]
  wire  writeMiss_st1 = cacheMiss_st1 & coreReq_st1_isWrite; // @[DCache.scala 156:37]
  wire  writeHitSubWord_st1 = writeHit_st1 & byteEn_st1; // @[DCache.scala 157:42]
  reg  writeMiss_st2; // @[DCache.scala 160:30]
  reg  writeMissSubWord_st2; // @[DCache.scala 161:37]
  reg  writeMiss_st3; // @[DCache.scala 162:30]
  reg  readHit_st2; // @[DCache.scala 164:28]
  reg  readHit_st2_REG; // @[DCache.scala 165:56]
  reg  readHit_st3; // @[DCache.scala 167:28]
  reg  writeHit_st2; // @[DCache.scala 168:29]
  reg  writeHit_st3; // @[DCache.scala 169:29]
  reg  bankConflict_st2; // @[DCache.scala 171:33]
  reg [7:0] arbDataCrsbarSel1H_st2_0; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_1; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_2; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_3; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_4; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_5; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_6; // @[DCache.scala 172:39]
  reg [7:0] arbDataCrsbarSel1H_st2_7; // @[DCache.scala 172:39]
  reg [3:0] arbAddrCrsbarOut_st2_0_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_1_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_2_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_3_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_4_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_5_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_6_wordOffset1H; // @[DCache.scala 173:37]
  reg [3:0] arbAddrCrsbarOut_st2_7_wordOffset1H; // @[DCache.scala 173:37]
  reg  arbArrayEn_st2_0; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_1; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_2; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_3; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_4; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_5; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_6; // @[DCache.scala 174:31]
  reg  arbArrayEn_st2_7; // @[DCache.scala 174:31]
  reg [7:0] arbDataCrsbarSel1H_st3_0; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_1; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_2; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_3; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_4; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_5; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_6; // @[DCache.scala 176:39]
  reg [7:0] arbDataCrsbarSel1H_st3_7; // @[DCache.scala 176:39]
  wire  _memRsp_Q_io_deq_ready_T_1 = ~(readHit_st2 | writeHit_st2); // @[DCache.scala 180:61]
  wire  _T_2 = memRsp_Q_io_deq_ready & memRsp_Q_io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _T_4 = _T_2 | memRsp_Q_io_deq_valid & BankConfArb_io_bankConflict; // @[DCache.scala 188:85]
  reg [31:0] r_0_0; // @[Reg.scala 16:16]
  reg [31:0] r_0_1; // @[Reg.scala 16:16]
  reg [31:0] r_0_2; // @[Reg.scala 16:16]
  reg [31:0] r_0_3; // @[Reg.scala 16:16]
  reg [31:0] r_0_4; // @[Reg.scala 16:16]
  reg [31:0] r_0_5; // @[Reg.scala 16:16]
  reg [31:0] r_0_6; // @[Reg.scala 16:16]
  reg [31:0] r_0_7; // @[Reg.scala 16:16]
  wire [31:0] memRspData_st1_0_0 = memRsp_Q_io_deq_bits_d_data_0; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_1 = memRsp_Q_io_deq_bits_d_data_1; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_2 = memRsp_Q_io_deq_bits_d_data_2; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_3 = memRsp_Q_io_deq_bits_d_data_3; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_4 = memRsp_Q_io_deq_bits_d_data_4; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_5 = memRsp_Q_io_deq_bits_d_data_5; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_6 = memRsp_Q_io_deq_bits_d_data_6; // @[DCache.scala 181:28 185:34]
  wire [31:0] memRspData_st1_0_7 = memRsp_Q_io_deq_bits_d_data_7; // @[DCache.scala 181:28 185:34]
  wire  _MshrAccess_io_missReq_valid_T_2 = _readHit_st1_T | coreReq_st1_isWrite & byteEn_st1; // @[DCache.scala 192:27]
  wire [15:0] MshrAccess_io_missReq_bits_targetInfo_lo_lo = {coreReq_st1_perLaneAddr_1_activeMask,
    coreReq_st1_perLaneAddr_1_blockOffset,4'hf,coreReq_st1_perLaneAddr_0_activeMask,
    coreReq_st1_perLaneAddr_0_blockOffset,4'hf}; // @[DCache.scala 199:64]
  wire [31:0] MshrAccess_io_missReq_bits_targetInfo_lo = {coreReq_st1_perLaneAddr_3_activeMask,
    coreReq_st1_perLaneAddr_3_blockOffset,4'hf,coreReq_st1_perLaneAddr_2_activeMask,
    coreReq_st1_perLaneAddr_2_blockOffset,4'hf,MshrAccess_io_missReq_bits_targetInfo_lo_lo}; // @[DCache.scala 199:64]
  wire [15:0] MshrAccess_io_missReq_bits_targetInfo_hi_lo = {coreReq_st1_perLaneAddr_5_activeMask,
    coreReq_st1_perLaneAddr_5_blockOffset,4'hf,coreReq_st1_perLaneAddr_4_activeMask,
    coreReq_st1_perLaneAddr_4_blockOffset,4'hf}; // @[DCache.scala 199:64]
  wire [32:0] MshrAccess_io_missReq_bits_targetInfo_hi = {coreReq_st1_isWrite,coreReq_st1_perLaneAddr_7_activeMask,
    coreReq_st1_perLaneAddr_7_blockOffset,4'hf,coreReq_st1_perLaneAddr_6_activeMask,
    coreReq_st1_perLaneAddr_6_blockOffset,4'hf,MshrAccess_io_missReq_bits_targetInfo_hi_lo}; // @[DCache.scala 199:64]
  reg  missRspTILaneMask_st2_0; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_1; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_2; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_3; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_4; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_5; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_6; // @[DCache.scala 207:38]
  reg  missRspTILaneMask_st2_7; // @[DCache.scala 207:38]
  reg [1:0] memRspInstrId_st2; // @[DCache.scala 208:34]
  reg  readMissRspCnter; // @[DCache.scala 210:91]
  wire  _MshrAccess_io_missRspOut_ready_T = ~missRspTI_st1_isWrite; // @[DCache.scala 213:6]
  wire [2:0] _coreRsp_QAlmstFull_T_1 = 3'h4 - 3'h2; // @[DCache.scala 332:73]
  wire  coreRsp_QAlmstFull = coreRsp_Q_io_count == _coreRsp_QAlmstFull_T_1; // @[DCache.scala 332:44]
  wire  _MshrAccess_io_missRspOut_ready_T_4 = ~missRspTI_st1_isWrite & ~BankConfArb_io_bankConflict & ~
    coreRsp_QAlmstFull; // @[DCache.scala 213:60]
  wire  _MshrAccess_io_missRspOut_ready_T_7 = missRspTI_st1_isWrite & ~WriteDataBuf_io_wdbAlmostFull; // @[DCache.scala 216:28]
  wire  _readMissRsp_st1_T = MshrAccess_io_missRspOut_ready & MshrAccess_io_missRspOut_valid; // @[Decoupled.scala 50:35]
  reg  readMissRsp_st2; // @[DCache.scala 223:32]
  reg  writeMissRsp_st2; // @[DCache.scala 224:33]
  wire  _T_5 = ~readMissRspCnter; // @[DCache.scala 225:25]
  reg  REG; // @[DCache.scala 226:16]
  reg [26:0] REG_1; // @[DCache.scala 227:13]
  wire  _T_8 = REG_1 != MshrAccess_io_missRspOut_bits_blockAddr; // @[DCache.scala 227:29]
  wire  _T_9 = ~REG & missRspFromMshr_st1 | _T_8; // @[DCache.scala 226:62]
  wire  _T_10 = _T_9 & missRspFromMshr_st1; // @[DCache.scala 227:49]
  wire  _T_11 = ~readMissRspCnter & _T_10; // @[DCache.scala 225:50]
  reg  missRspWriteEnable_REG; // @[DCache.scala 232:36]
  reg [26:0] missRspWriteEnable_REG_1; // @[DCache.scala 233:13]
  wire  _missRspWriteEnable_T_2 = missRspWriteEnable_REG_1 != MshrAccess_io_missRspOut_bits_blockAddr; // @[DCache.scala 233:29]
  wire  _missRspWriteEnable_T_3 = ~missRspWriteEnable_REG & missRspFromMshr_st1 | _missRspWriteEnable_T_2; // @[DCache.scala 232:82]
  wire  missRspWriteEnable = _missRspWriteEnable_T_3 & missRspFromMshr_st1 | _T_5; // @[DCache.scala 233:73]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T = writeHit_st2 & arbArrayEn_st2_0; // @[DCache.scala 249:20]
  wire [31:0] _DataAccessesRRsp_T__0 = missRspWriteEnable ? memRspData_st1_0_0 : DataCorssBar_io_DataOut_0; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__1 = missRspWriteEnable ? memRspData_st1_0_1 : DataCorssBar_io_DataOut_1; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__2 = missRspWriteEnable ? memRspData_st1_0_2 : DataCorssBar_io_DataOut_2; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__3 = missRspWriteEnable ? memRspData_st1_0_3 : DataCorssBar_io_DataOut_3; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__4 = missRspWriteEnable ? memRspData_st1_0_4 : DataCorssBar_io_DataOut_4; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__5 = missRspWriteEnable ? memRspData_st1_0_5 : DataCorssBar_io_DataOut_5; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__6 = missRspWriteEnable ? memRspData_st1_0_6 : DataCorssBar_io_DataOut_6; // @[DCache.scala 255:35]
  wire [31:0] _DataAccessesRRsp_T__7 = missRspWriteEnable ? memRspData_st1_0_7 : DataCorssBar_io_DataOut_7; // @[DCache.scala 255:35]
  wire [5:0] DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 = {memRsp_Q_io_deq_bits_d_addr[9:5],wayIdxReplace_st0}; // @[Cat.scala 31:58]
  wire [5:0] DataAccessesRRsp_DAWtSetIdxWtHitCase_st2 = {coreReq_st2_setIdx,wayIdxAtHit_st2}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_2 = writeHitSubWord_st1 & writeSubWordBank_st1[0]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_0 = {DataAccessesRRsp_DataAccess_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_io_r_resp_data_2,DataAccessesRRsp_DataAccess_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_2 = writeHit_st2 & arbArrayEn_st2_1; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_6 = writeHitSubWord_st1 & writeSubWordBank_st1[1]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_1 = {DataAccessesRRsp_DataAccess_1_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_1_io_r_resp_data_2,DataAccessesRRsp_DataAccess_1_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_1_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_4 = writeHit_st2 & arbArrayEn_st2_2; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_10 = writeHitSubWord_st1 & writeSubWordBank_st1[2]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_2 = {DataAccessesRRsp_DataAccess_2_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_2_io_r_resp_data_2,DataAccessesRRsp_DataAccess_2_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_2_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_6 = writeHit_st2 & arbArrayEn_st2_3; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_14 = writeHitSubWord_st1 & writeSubWordBank_st1[3]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_3 = {DataAccessesRRsp_DataAccess_3_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_3_io_r_resp_data_2,DataAccessesRRsp_DataAccess_3_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_3_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_8 = writeHit_st2 & arbArrayEn_st2_4; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_18 = writeHitSubWord_st1 & writeSubWordBank_st1[4]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_4 = {DataAccessesRRsp_DataAccess_4_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_4_io_r_resp_data_2,DataAccessesRRsp_DataAccess_4_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_4_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_10 = writeHit_st2 & arbArrayEn_st2_5; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_22 = writeHitSubWord_st1 & writeSubWordBank_st1[5]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_5 = {DataAccessesRRsp_DataAccess_5_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_5_io_r_resp_data_2,DataAccessesRRsp_DataAccess_5_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_5_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_12 = writeHit_st2 & arbArrayEn_st2_6; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_26 = writeHitSubWord_st1 & writeSubWordBank_st1[6]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_6 = {DataAccessesRRsp_DataAccess_6_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_6_io_r_resp_data_2,DataAccessesRRsp_DataAccess_6_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_6_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire  _DataAccessesRRsp_DataAccess_io_w_req_valid_T_14 = writeHit_st2 & arbArrayEn_st2_7; // @[DCache.scala 249:20]
  wire  _DataAccessesRRsp_DataAccess_io_r_req_valid_T_30 = writeHitSubWord_st1 & writeSubWordBank_st1[7]; // @[DCache.scala 286:28]
  wire [31:0] DataAccessesRRsp_7 = {DataAccessesRRsp_DataAccess_7_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_7_io_r_resp_data_2,DataAccessesRRsp_DataAccess_7_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_7_io_r_resp_data_0}; // @[Cat.scala 31:58]
  reg [31:0] dataAccess_data_st3_0; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_1; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_2; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_3; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_4; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_5; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_6; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st3_7; // @[Reg.scala 16:16]
  wire [31:0] _T_14_0 = coreReq_st2_isWrite ? coreReq_st2_data_0 : dataAccess_data_st3_0; // @[DCache.scala 303:8]
  wire [31:0] _T_14_1 = coreReq_st2_isWrite ? coreReq_st2_data_1 : dataAccess_data_st3_1; // @[DCache.scala 303:8]
  wire [31:0] _T_14_2 = coreReq_st2_isWrite ? coreReq_st2_data_2 : dataAccess_data_st3_2; // @[DCache.scala 303:8]
  wire [31:0] _T_14_3 = coreReq_st2_isWrite ? coreReq_st2_data_3 : dataAccess_data_st3_3; // @[DCache.scala 303:8]
  wire [31:0] _T_14_4 = coreReq_st2_isWrite ? coreReq_st2_data_4 : dataAccess_data_st3_4; // @[DCache.scala 303:8]
  wire [31:0] _T_14_5 = coreReq_st2_isWrite ? coreReq_st2_data_5 : dataAccess_data_st3_5; // @[DCache.scala 303:8]
  wire [31:0] _T_14_6 = coreReq_st2_isWrite ? coreReq_st2_data_6 : dataAccess_data_st3_6; // @[DCache.scala 303:8]
  wire [31:0] _T_14_7 = coreReq_st2_isWrite ? coreReq_st2_data_7 : dataAccess_data_st3_7; // @[DCache.scala 303:8]
  wire  _io_coreReq_ready_T_2 = ~missRspFromMshr_st1; // @[DCache.scala 337:5]
  wire  _io_coreReq_ready_T_3 = ~(BankConfArb_io_bankConflict & readHit_st1) & _io_coreReq_ready_T_2; // @[DCache.scala 336:68]
  wire  _io_coreReq_ready_T_7 = ~(readHit_st1 & coreRsp_QAlmstFull); // @[DCache.scala 338:5]
  wire  _io_coreReq_ready_T_8 = _io_coreReq_ready_T_3 & ~io_memRsp_valid & _io_coreReq_ready_T_7; // @[DCache.scala 337:45]
  wire  _io_coreReq_ready_T_10 = ~(coreReq_st1_isWrite & WriteDataBuf_io_wdbAlmostFull); // @[DCache.scala 339:5]
  wire  _io_coreReq_ready_T_11 = _io_coreReq_ready_T_8 & _io_coreReq_ready_T_10; // @[DCache.scala 338:41]
  wire  _io_coreReq_ready_T_13 = ~(readHit_st2 & coreReq_st1_isWrite); // @[DCache.scala 340:5]
  wire  _io_coreReq_ready_T_14 = _io_coreReq_ready_T_11 & _io_coreReq_ready_T_13; // @[DCache.scala 339:60]
  wire  _WriteDataBuf_io_inputBus_valid_T_1 = writeMissRsp_st2 & missRspTI_st1_isWrite; // @[DCache.scala 345:23]
  wire [255:0] _T_19 = {DataCorssBar_io_DataOut_7,DataCorssBar_io_DataOut_6,DataCorssBar_io_DataOut_5,
    DataCorssBar_io_DataOut_4,DataCorssBar_io_DataOut_3,DataCorssBar_io_DataOut_2,DataCorssBar_io_DataOut_1,
    DataCorssBar_io_DataOut_0}; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_0_0 = _T_19[7:0]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_0_1 = _T_19[15:8]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_0_2 = _T_19[23:16]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_0_3 = _T_19[31:24]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_1_0 = _T_19[39:32]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_1_1 = _T_19[47:40]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_1_2 = _T_19[55:48]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_1_3 = _T_19[63:56]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_2_0 = _T_19[71:64]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_2_1 = _T_19[79:72]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_2_2 = _T_19[87:80]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_2_3 = _T_19[95:88]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_3_0 = _T_19[103:96]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_3_1 = _T_19[111:104]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_3_2 = _T_19[119:112]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_3_3 = _T_19[127:120]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_4_0 = _T_19[135:128]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_4_1 = _T_19[143:136]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_4_2 = _T_19[151:144]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_4_3 = _T_19[159:152]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_5_0 = _T_19[167:160]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_5_1 = _T_19[175:168]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_5_2 = _T_19[183:176]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_5_3 = _T_19[191:184]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_6_0 = _T_19[199:192]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_6_1 = _T_19[207:200]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_6_2 = _T_19[215:208]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_6_3 = _T_19[223:216]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_7_0 = _T_19[231:224]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_7_1 = _T_19[239:232]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_7_2 = _T_19[247:240]; // @[DCache.scala 347:58]
  wire [7:0] DataCrsbarToWdb_st2_7_3 = _T_19[255:248]; // @[DCache.scala 347:58]
  wire [3:0] perWordByteMask_0 = arbArrayEn_st2_0 ? arbAddrCrsbarOut_st2_0_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_0_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_0_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_0_0_T_3 = perWordByteMask_0[0] ? DataCrsbarToWdb_st2_0_0 : {{7'd0},
    DataAccessesRRsp_0[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_0_1_T_3 = perWordByteMask_0[1] ? DataCrsbarToWdb_st2_0_1 : {{7'd0},
    DataAccessesRRsp_0[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_0_2_T_3 = perWordByteMask_0[2] ? DataCrsbarToWdb_st2_0_2 : {{7'd0},
    DataAccessesRRsp_0[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_0_3_T_3 = perWordByteMask_0[3] ? DataCrsbarToWdb_st2_0_3 : {{7'd0},
    DataAccessesRRsp_0[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_1 = arbArrayEn_st2_1 ? arbAddrCrsbarOut_st2_1_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_1_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_1_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_1_0_T_3 = perWordByteMask_1[0] ? DataCrsbarToWdb_st2_1_0 : {{7'd0},
    DataAccessesRRsp_1[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_1_1_T_3 = perWordByteMask_1[1] ? DataCrsbarToWdb_st2_1_1 : {{7'd0},
    DataAccessesRRsp_1[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_1_2_T_3 = perWordByteMask_1[2] ? DataCrsbarToWdb_st2_1_2 : {{7'd0},
    DataAccessesRRsp_1[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_1_3_T_3 = perWordByteMask_1[3] ? DataCrsbarToWdb_st2_1_3 : {{7'd0},
    DataAccessesRRsp_1[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_2 = arbArrayEn_st2_2 ? arbAddrCrsbarOut_st2_2_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_2_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_2_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_2_0_T_3 = perWordByteMask_2[0] ? DataCrsbarToWdb_st2_2_0 : {{7'd0},
    DataAccessesRRsp_2[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_2_1_T_3 = perWordByteMask_2[1] ? DataCrsbarToWdb_st2_2_1 : {{7'd0},
    DataAccessesRRsp_2[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_2_2_T_3 = perWordByteMask_2[2] ? DataCrsbarToWdb_st2_2_2 : {{7'd0},
    DataAccessesRRsp_2[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_2_3_T_3 = perWordByteMask_2[3] ? DataCrsbarToWdb_st2_2_3 : {{7'd0},
    DataAccessesRRsp_2[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_3 = arbArrayEn_st2_3 ? arbAddrCrsbarOut_st2_3_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_3_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_3_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_3_0_T_3 = perWordByteMask_3[0] ? DataCrsbarToWdb_st2_3_0 : {{7'd0},
    DataAccessesRRsp_3[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_3_1_T_3 = perWordByteMask_3[1] ? DataCrsbarToWdb_st2_3_1 : {{7'd0},
    DataAccessesRRsp_3[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_3_2_T_3 = perWordByteMask_3[2] ? DataCrsbarToWdb_st2_3_2 : {{7'd0},
    DataAccessesRRsp_3[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_3_3_T_3 = perWordByteMask_3[3] ? DataCrsbarToWdb_st2_3_3 : {{7'd0},
    DataAccessesRRsp_3[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_4 = arbArrayEn_st2_4 ? arbAddrCrsbarOut_st2_4_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_4_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_4_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_4_0_T_3 = perWordByteMask_4[0] ? DataCrsbarToWdb_st2_4_0 : {{7'd0},
    DataAccessesRRsp_4[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_4_1_T_3 = perWordByteMask_4[1] ? DataCrsbarToWdb_st2_4_1 : {{7'd0},
    DataAccessesRRsp_4[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_4_2_T_3 = perWordByteMask_4[2] ? DataCrsbarToWdb_st2_4_2 : {{7'd0},
    DataAccessesRRsp_4[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_4_3_T_3 = perWordByteMask_4[3] ? DataCrsbarToWdb_st2_4_3 : {{7'd0},
    DataAccessesRRsp_4[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_5 = arbArrayEn_st2_5 ? arbAddrCrsbarOut_st2_5_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_5_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_5_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_5_0_T_3 = perWordByteMask_5[0] ? DataCrsbarToWdb_st2_5_0 : {{7'd0},
    DataAccessesRRsp_5[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_5_1_T_3 = perWordByteMask_5[1] ? DataCrsbarToWdb_st2_5_1 : {{7'd0},
    DataAccessesRRsp_5[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_5_2_T_3 = perWordByteMask_5[2] ? DataCrsbarToWdb_st2_5_2 : {{7'd0},
    DataAccessesRRsp_5[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_5_3_T_3 = perWordByteMask_5[3] ? DataCrsbarToWdb_st2_5_3 : {{7'd0},
    DataAccessesRRsp_5[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_6 = arbArrayEn_st2_6 ? arbAddrCrsbarOut_st2_6_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_6_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_6_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_6_0_T_3 = perWordByteMask_6[0] ? DataCrsbarToWdb_st2_6_0 : {{7'd0},
    DataAccessesRRsp_6[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_6_1_T_3 = perWordByteMask_6[1] ? DataCrsbarToWdb_st2_6_1 : {{7'd0},
    DataAccessesRRsp_6[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_6_2_T_3 = perWordByteMask_6[2] ? DataCrsbarToWdb_st2_6_2 : {{7'd0},
    DataAccessesRRsp_6[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_6_3_T_3 = perWordByteMask_6[3] ? DataCrsbarToWdb_st2_6_3 : {{7'd0},
    DataAccessesRRsp_6[3]}; // @[DCache.scala 367:18]
  wire [3:0] perWordByteMask_7 = arbArrayEn_st2_7 ? arbAddrCrsbarOut_st2_7_wordOffset1H : 4'h0; // @[DCache.scala 352:12]
  wire [3:0] _WriteDataBuf_io_inputBus_bits_mask_7_T_2 = writeMissSubWord_st2 ? arbAddrCrsbarOut_st2_7_wordOffset1H : 4'hf
    ; // @[DCache.scala 360:16]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_7_0_T_3 = perWordByteMask_7[0] ? DataCrsbarToWdb_st2_7_0 : {{7'd0},
    DataAccessesRRsp_7[0]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_7_1_T_3 = perWordByteMask_7[1] ? DataCrsbarToWdb_st2_7_1 : {{7'd0},
    DataAccessesRRsp_7[1]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_7_2_T_3 = perWordByteMask_7[2] ? DataCrsbarToWdb_st2_7_2 : {{7'd0},
    DataAccessesRRsp_7[2]}; // @[DCache.scala 367:18]
  wire [7:0] _WriteDataBuf_io_inputBus_bits_data_7_3_T_3 = perWordByteMask_7[3] ? DataCrsbarToWdb_st2_7_3 : {{7'd0},
    DataAccessesRRsp_7[3]}; // @[DCache.scala 367:18]
  wire [26:0] WriteDataBuf_io_inputBus_bits_addr_hi = {coreReq_st2_tag,coreReq_st2_setIdx}; // @[Cat.scala 31:58]
  wire [7:0] _wdbMemReq_a_opcode_T = {WriteDataBuf_io_outputBus_bits_mask_0,WriteDataBuf_io_outputBus_bits_mask_1,
    WriteDataBuf_io_outputBus_bits_mask_2,WriteDataBuf_io_outputBus_bits_mask_3,WriteDataBuf_io_outputBus_bits_mask_4,
    WriteDataBuf_io_outputBus_bits_mask_5,WriteDataBuf_io_outputBus_bits_mask_6,WriteDataBuf_io_outputBus_bits_mask_7}; // @[Cat.scala 31:58]
  wire [63:0] lo_lo_1 = {WriteDataBuf_io_outputBus_bits_data_1_3,WriteDataBuf_io_outputBus_bits_data_1_2,
    WriteDataBuf_io_outputBus_bits_data_1_1,WriteDataBuf_io_outputBus_bits_data_1_0,
    WriteDataBuf_io_outputBus_bits_data_0_3,WriteDataBuf_io_outputBus_bits_data_0_2,
    WriteDataBuf_io_outputBus_bits_data_0_1,WriteDataBuf_io_outputBus_bits_data_0_0}; // @[DCache.scala 396:48]
  wire [127:0] lo_1 = {WriteDataBuf_io_outputBus_bits_data_3_3,WriteDataBuf_io_outputBus_bits_data_3_2,
    WriteDataBuf_io_outputBus_bits_data_3_1,WriteDataBuf_io_outputBus_bits_data_3_0,
    WriteDataBuf_io_outputBus_bits_data_2_3,WriteDataBuf_io_outputBus_bits_data_2_2,
    WriteDataBuf_io_outputBus_bits_data_2_1,WriteDataBuf_io_outputBus_bits_data_2_0,lo_lo_1}; // @[DCache.scala 396:48]
  wire [63:0] hi_lo_1 = {WriteDataBuf_io_outputBus_bits_data_5_3,WriteDataBuf_io_outputBus_bits_data_5_2,
    WriteDataBuf_io_outputBus_bits_data_5_1,WriteDataBuf_io_outputBus_bits_data_5_0,
    WriteDataBuf_io_outputBus_bits_data_4_3,WriteDataBuf_io_outputBus_bits_data_4_2,
    WriteDataBuf_io_outputBus_bits_data_4_1,WriteDataBuf_io_outputBus_bits_data_4_0}; // @[DCache.scala 396:48]
  wire [255:0] _T_52 = {WriteDataBuf_io_outputBus_bits_data_7_3,WriteDataBuf_io_outputBus_bits_data_7_2,
    WriteDataBuf_io_outputBus_bits_data_7_1,WriteDataBuf_io_outputBus_bits_data_7_0,
    WriteDataBuf_io_outputBus_bits_data_6_3,WriteDataBuf_io_outputBus_bits_data_6_2,
    WriteDataBuf_io_outputBus_bits_data_6_1,WriteDataBuf_io_outputBus_bits_data_6_0,hi_lo_1,lo_1}; // @[DCache.scala 396:48]
  BankConflictArbiter BankConfArb ( // @[DCache.scala 85:27]
    .clock(BankConfArb_clock),
    .reset(BankConfArb_reset),
    .io_coreReqArb_isWrite(BankConfArb_io_coreReqArb_isWrite),
    .io_coreReqArb_enable(BankConfArb_io_coreReqArb_enable),
    .io_coreReqArb_perLaneAddr_0_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_0_activeMask),
    .io_coreReqArb_perLaneAddr_0_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_0_blockOffset),
    .io_coreReqArb_perLaneAddr_0_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_0_wordOffset1H),
    .io_coreReqArb_perLaneAddr_1_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_1_activeMask),
    .io_coreReqArb_perLaneAddr_1_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_1_blockOffset),
    .io_coreReqArb_perLaneAddr_1_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_1_wordOffset1H),
    .io_coreReqArb_perLaneAddr_2_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_2_activeMask),
    .io_coreReqArb_perLaneAddr_2_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_2_blockOffset),
    .io_coreReqArb_perLaneAddr_2_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_2_wordOffset1H),
    .io_coreReqArb_perLaneAddr_3_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_3_activeMask),
    .io_coreReqArb_perLaneAddr_3_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_3_blockOffset),
    .io_coreReqArb_perLaneAddr_3_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_3_wordOffset1H),
    .io_coreReqArb_perLaneAddr_4_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_4_activeMask),
    .io_coreReqArb_perLaneAddr_4_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_4_blockOffset),
    .io_coreReqArb_perLaneAddr_4_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_4_wordOffset1H),
    .io_coreReqArb_perLaneAddr_5_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_5_activeMask),
    .io_coreReqArb_perLaneAddr_5_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_5_blockOffset),
    .io_coreReqArb_perLaneAddr_5_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_5_wordOffset1H),
    .io_coreReqArb_perLaneAddr_6_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_6_activeMask),
    .io_coreReqArb_perLaneAddr_6_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_6_blockOffset),
    .io_coreReqArb_perLaneAddr_6_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_6_wordOffset1H),
    .io_coreReqArb_perLaneAddr_7_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_7_activeMask),
    .io_coreReqArb_perLaneAddr_7_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_7_blockOffset),
    .io_coreReqArb_perLaneAddr_7_wordOffset1H(BankConfArb_io_coreReqArb_perLaneAddr_7_wordOffset1H),
    .io_dataCrsbarSel1H_0(BankConfArb_io_dataCrsbarSel1H_0),
    .io_dataCrsbarSel1H_1(BankConfArb_io_dataCrsbarSel1H_1),
    .io_dataCrsbarSel1H_2(BankConfArb_io_dataCrsbarSel1H_2),
    .io_dataCrsbarSel1H_3(BankConfArb_io_dataCrsbarSel1H_3),
    .io_dataCrsbarSel1H_4(BankConfArb_io_dataCrsbarSel1H_4),
    .io_dataCrsbarSel1H_5(BankConfArb_io_dataCrsbarSel1H_5),
    .io_dataCrsbarSel1H_6(BankConfArb_io_dataCrsbarSel1H_6),
    .io_dataCrsbarSel1H_7(BankConfArb_io_dataCrsbarSel1H_7),
    .io_addrCrsbarOut_0_wordOffset1H(BankConfArb_io_addrCrsbarOut_0_wordOffset1H),
    .io_addrCrsbarOut_1_wordOffset1H(BankConfArb_io_addrCrsbarOut_1_wordOffset1H),
    .io_addrCrsbarOut_2_wordOffset1H(BankConfArb_io_addrCrsbarOut_2_wordOffset1H),
    .io_addrCrsbarOut_3_wordOffset1H(BankConfArb_io_addrCrsbarOut_3_wordOffset1H),
    .io_addrCrsbarOut_4_wordOffset1H(BankConfArb_io_addrCrsbarOut_4_wordOffset1H),
    .io_addrCrsbarOut_5_wordOffset1H(BankConfArb_io_addrCrsbarOut_5_wordOffset1H),
    .io_addrCrsbarOut_6_wordOffset1H(BankConfArb_io_addrCrsbarOut_6_wordOffset1H),
    .io_addrCrsbarOut_7_wordOffset1H(BankConfArb_io_addrCrsbarOut_7_wordOffset1H),
    .io_dataArrayEn_0(BankConfArb_io_dataArrayEn_0),
    .io_dataArrayEn_1(BankConfArb_io_dataArrayEn_1),
    .io_dataArrayEn_2(BankConfArb_io_dataArrayEn_2),
    .io_dataArrayEn_3(BankConfArb_io_dataArrayEn_3),
    .io_dataArrayEn_4(BankConfArb_io_dataArrayEn_4),
    .io_dataArrayEn_5(BankConfArb_io_dataArrayEn_5),
    .io_dataArrayEn_6(BankConfArb_io_dataArrayEn_6),
    .io_dataArrayEn_7(BankConfArb_io_dataArrayEn_7),
    .io_activeLane_0(BankConfArb_io_activeLane_0),
    .io_activeLane_1(BankConfArb_io_activeLane_1),
    .io_activeLane_2(BankConfArb_io_activeLane_2),
    .io_activeLane_3(BankConfArb_io_activeLane_3),
    .io_activeLane_4(BankConfArb_io_activeLane_4),
    .io_activeLane_5(BankConfArb_io_activeLane_5),
    .io_activeLane_6(BankConfArb_io_activeLane_6),
    .io_activeLane_7(BankConfArb_io_activeLane_7),
    .io_bankConflict(BankConfArb_io_bankConflict)
  );
  MSHR_1 MshrAccess ( // @[DCache.scala 87:26]
    .clock(MshrAccess_clock),
    .reset(MshrAccess_reset),
    .io_missReq_ready(MshrAccess_io_missReq_ready),
    .io_missReq_valid(MshrAccess_io_missReq_valid),
    .io_missReq_bits_blockAddr(MshrAccess_io_missReq_bits_blockAddr),
    .io_missReq_bits_instrId(MshrAccess_io_missReq_bits_instrId),
    .io_missReq_bits_targetInfo(MshrAccess_io_missReq_bits_targetInfo),
    .io_missRspIn_ready(MshrAccess_io_missRspIn_ready),
    .io_missRspIn_valid(MshrAccess_io_missRspIn_valid),
    .io_missRspIn_bits_blockAddr(MshrAccess_io_missRspIn_bits_blockAddr),
    .io_missRspOut_ready(MshrAccess_io_missRspOut_ready),
    .io_missRspOut_valid(MshrAccess_io_missRspOut_valid),
    .io_missRspOut_bits_targetInfo(MshrAccess_io_missRspOut_bits_targetInfo),
    .io_missRspOut_bits_blockAddr(MshrAccess_io_missRspOut_bits_blockAddr),
    .io_missRspOut_bits_instrId(MshrAccess_io_missRspOut_bits_instrId),
    .io_miss2mem_ready(MshrAccess_io_miss2mem_ready),
    .io_miss2mem_valid(MshrAccess_io_miss2mem_valid),
    .io_miss2mem_bits_blockAddr(MshrAccess_io_miss2mem_bits_blockAddr),
    .io_miss2mem_bits_instrId(MshrAccess_io_miss2mem_bits_instrId)
  );
  L1TagAccess TagAccess ( // @[DCache.scala 90:25]
    .clock(TagAccess_clock),
    .reset(TagAccess_reset),
    .io_r_req_valid(TagAccess_io_r_req_valid),
    .io_r_req_bits_setIdx(TagAccess_io_r_req_bits_setIdx),
    .io_tagFromCore_st1(TagAccess_io_tagFromCore_st1),
    .io_coreReqReady(TagAccess_io_coreReqReady),
    .io_w_req_valid(TagAccess_io_w_req_valid),
    .io_w_req_bits_setIdx(TagAccess_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(TagAccess_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(TagAccess_io_w_req_bits_data_1),
    .io_waymaskReplacement(TagAccess_io_waymaskReplacement),
    .io_waymaskHit_st1(TagAccess_io_waymaskHit_st1),
    .io_hit_st1(TagAccess_io_hit_st1)
  );
  DataCrossbar DataCorssBar ( // @[DCache.scala 91:28]
    .io_DataIn_0(DataCorssBar_io_DataIn_0),
    .io_DataIn_1(DataCorssBar_io_DataIn_1),
    .io_DataIn_2(DataCorssBar_io_DataIn_2),
    .io_DataIn_3(DataCorssBar_io_DataIn_3),
    .io_DataIn_4(DataCorssBar_io_DataIn_4),
    .io_DataIn_5(DataCorssBar_io_DataIn_5),
    .io_DataIn_6(DataCorssBar_io_DataIn_6),
    .io_DataIn_7(DataCorssBar_io_DataIn_7),
    .io_DataOut_0(DataCorssBar_io_DataOut_0),
    .io_DataOut_1(DataCorssBar_io_DataOut_1),
    .io_DataOut_2(DataCorssBar_io_DataOut_2),
    .io_DataOut_3(DataCorssBar_io_DataOut_3),
    .io_DataOut_4(DataCorssBar_io_DataOut_4),
    .io_DataOut_5(DataCorssBar_io_DataOut_5),
    .io_DataOut_6(DataCorssBar_io_DataOut_6),
    .io_DataOut_7(DataCorssBar_io_DataOut_7),
    .io_Select1H_0(DataCorssBar_io_Select1H_0),
    .io_Select1H_1(DataCorssBar_io_Select1H_1),
    .io_Select1H_2(DataCorssBar_io_Select1H_2),
    .io_Select1H_3(DataCorssBar_io_Select1H_3),
    .io_Select1H_4(DataCorssBar_io_Select1H_4),
    .io_Select1H_5(DataCorssBar_io_Select1H_5),
    .io_Select1H_6(DataCorssBar_io_Select1H_6),
    .io_Select1H_7(DataCorssBar_io_Select1H_7)
  );
  WDB WriteDataBuf ( // @[DCache.scala 92:28]
    .clock(WriteDataBuf_clock),
    .reset(WriteDataBuf_reset),
    .io_inputBus_ready(WriteDataBuf_io_inputBus_ready),
    .io_inputBus_valid(WriteDataBuf_io_inputBus_valid),
    .io_inputBus_bits_mask_0(WriteDataBuf_io_inputBus_bits_mask_0),
    .io_inputBus_bits_mask_1(WriteDataBuf_io_inputBus_bits_mask_1),
    .io_inputBus_bits_mask_2(WriteDataBuf_io_inputBus_bits_mask_2),
    .io_inputBus_bits_mask_3(WriteDataBuf_io_inputBus_bits_mask_3),
    .io_inputBus_bits_mask_4(WriteDataBuf_io_inputBus_bits_mask_4),
    .io_inputBus_bits_mask_5(WriteDataBuf_io_inputBus_bits_mask_5),
    .io_inputBus_bits_mask_6(WriteDataBuf_io_inputBus_bits_mask_6),
    .io_inputBus_bits_mask_7(WriteDataBuf_io_inputBus_bits_mask_7),
    .io_inputBus_bits_addr(WriteDataBuf_io_inputBus_bits_addr),
    .io_inputBus_bits_data_0_0(WriteDataBuf_io_inputBus_bits_data_0_0),
    .io_inputBus_bits_data_0_1(WriteDataBuf_io_inputBus_bits_data_0_1),
    .io_inputBus_bits_data_0_2(WriteDataBuf_io_inputBus_bits_data_0_2),
    .io_inputBus_bits_data_0_3(WriteDataBuf_io_inputBus_bits_data_0_3),
    .io_inputBus_bits_data_1_0(WriteDataBuf_io_inputBus_bits_data_1_0),
    .io_inputBus_bits_data_1_1(WriteDataBuf_io_inputBus_bits_data_1_1),
    .io_inputBus_bits_data_1_2(WriteDataBuf_io_inputBus_bits_data_1_2),
    .io_inputBus_bits_data_1_3(WriteDataBuf_io_inputBus_bits_data_1_3),
    .io_inputBus_bits_data_2_0(WriteDataBuf_io_inputBus_bits_data_2_0),
    .io_inputBus_bits_data_2_1(WriteDataBuf_io_inputBus_bits_data_2_1),
    .io_inputBus_bits_data_2_2(WriteDataBuf_io_inputBus_bits_data_2_2),
    .io_inputBus_bits_data_2_3(WriteDataBuf_io_inputBus_bits_data_2_3),
    .io_inputBus_bits_data_3_0(WriteDataBuf_io_inputBus_bits_data_3_0),
    .io_inputBus_bits_data_3_1(WriteDataBuf_io_inputBus_bits_data_3_1),
    .io_inputBus_bits_data_3_2(WriteDataBuf_io_inputBus_bits_data_3_2),
    .io_inputBus_bits_data_3_3(WriteDataBuf_io_inputBus_bits_data_3_3),
    .io_inputBus_bits_data_4_0(WriteDataBuf_io_inputBus_bits_data_4_0),
    .io_inputBus_bits_data_4_1(WriteDataBuf_io_inputBus_bits_data_4_1),
    .io_inputBus_bits_data_4_2(WriteDataBuf_io_inputBus_bits_data_4_2),
    .io_inputBus_bits_data_4_3(WriteDataBuf_io_inputBus_bits_data_4_3),
    .io_inputBus_bits_data_5_0(WriteDataBuf_io_inputBus_bits_data_5_0),
    .io_inputBus_bits_data_5_1(WriteDataBuf_io_inputBus_bits_data_5_1),
    .io_inputBus_bits_data_5_2(WriteDataBuf_io_inputBus_bits_data_5_2),
    .io_inputBus_bits_data_5_3(WriteDataBuf_io_inputBus_bits_data_5_3),
    .io_inputBus_bits_data_6_0(WriteDataBuf_io_inputBus_bits_data_6_0),
    .io_inputBus_bits_data_6_1(WriteDataBuf_io_inputBus_bits_data_6_1),
    .io_inputBus_bits_data_6_2(WriteDataBuf_io_inputBus_bits_data_6_2),
    .io_inputBus_bits_data_6_3(WriteDataBuf_io_inputBus_bits_data_6_3),
    .io_inputBus_bits_data_7_0(WriteDataBuf_io_inputBus_bits_data_7_0),
    .io_inputBus_bits_data_7_1(WriteDataBuf_io_inputBus_bits_data_7_1),
    .io_inputBus_bits_data_7_2(WriteDataBuf_io_inputBus_bits_data_7_2),
    .io_inputBus_bits_data_7_3(WriteDataBuf_io_inputBus_bits_data_7_3),
    .io_inputBus_bits_instrId(WriteDataBuf_io_inputBus_bits_instrId),
    .io_inputBus_bits_bankConflict(WriteDataBuf_io_inputBus_bits_bankConflict),
    .io_inputBus_bits_subWordMissReq(WriteDataBuf_io_inputBus_bits_subWordMissReq),
    .io_inputBus_bits_subWordMissRsp(WriteDataBuf_io_inputBus_bits_subWordMissRsp),
    .io_outputBus_ready(WriteDataBuf_io_outputBus_ready),
    .io_outputBus_valid(WriteDataBuf_io_outputBus_valid),
    .io_outputBus_bits_mask_0(WriteDataBuf_io_outputBus_bits_mask_0),
    .io_outputBus_bits_mask_1(WriteDataBuf_io_outputBus_bits_mask_1),
    .io_outputBus_bits_mask_2(WriteDataBuf_io_outputBus_bits_mask_2),
    .io_outputBus_bits_mask_3(WriteDataBuf_io_outputBus_bits_mask_3),
    .io_outputBus_bits_mask_4(WriteDataBuf_io_outputBus_bits_mask_4),
    .io_outputBus_bits_mask_5(WriteDataBuf_io_outputBus_bits_mask_5),
    .io_outputBus_bits_mask_6(WriteDataBuf_io_outputBus_bits_mask_6),
    .io_outputBus_bits_mask_7(WriteDataBuf_io_outputBus_bits_mask_7),
    .io_outputBus_bits_addr(WriteDataBuf_io_outputBus_bits_addr),
    .io_outputBus_bits_data_0_0(WriteDataBuf_io_outputBus_bits_data_0_0),
    .io_outputBus_bits_data_0_1(WriteDataBuf_io_outputBus_bits_data_0_1),
    .io_outputBus_bits_data_0_2(WriteDataBuf_io_outputBus_bits_data_0_2),
    .io_outputBus_bits_data_0_3(WriteDataBuf_io_outputBus_bits_data_0_3),
    .io_outputBus_bits_data_1_0(WriteDataBuf_io_outputBus_bits_data_1_0),
    .io_outputBus_bits_data_1_1(WriteDataBuf_io_outputBus_bits_data_1_1),
    .io_outputBus_bits_data_1_2(WriteDataBuf_io_outputBus_bits_data_1_2),
    .io_outputBus_bits_data_1_3(WriteDataBuf_io_outputBus_bits_data_1_3),
    .io_outputBus_bits_data_2_0(WriteDataBuf_io_outputBus_bits_data_2_0),
    .io_outputBus_bits_data_2_1(WriteDataBuf_io_outputBus_bits_data_2_1),
    .io_outputBus_bits_data_2_2(WriteDataBuf_io_outputBus_bits_data_2_2),
    .io_outputBus_bits_data_2_3(WriteDataBuf_io_outputBus_bits_data_2_3),
    .io_outputBus_bits_data_3_0(WriteDataBuf_io_outputBus_bits_data_3_0),
    .io_outputBus_bits_data_3_1(WriteDataBuf_io_outputBus_bits_data_3_1),
    .io_outputBus_bits_data_3_2(WriteDataBuf_io_outputBus_bits_data_3_2),
    .io_outputBus_bits_data_3_3(WriteDataBuf_io_outputBus_bits_data_3_3),
    .io_outputBus_bits_data_4_0(WriteDataBuf_io_outputBus_bits_data_4_0),
    .io_outputBus_bits_data_4_1(WriteDataBuf_io_outputBus_bits_data_4_1),
    .io_outputBus_bits_data_4_2(WriteDataBuf_io_outputBus_bits_data_4_2),
    .io_outputBus_bits_data_4_3(WriteDataBuf_io_outputBus_bits_data_4_3),
    .io_outputBus_bits_data_5_0(WriteDataBuf_io_outputBus_bits_data_5_0),
    .io_outputBus_bits_data_5_1(WriteDataBuf_io_outputBus_bits_data_5_1),
    .io_outputBus_bits_data_5_2(WriteDataBuf_io_outputBus_bits_data_5_2),
    .io_outputBus_bits_data_5_3(WriteDataBuf_io_outputBus_bits_data_5_3),
    .io_outputBus_bits_data_6_0(WriteDataBuf_io_outputBus_bits_data_6_0),
    .io_outputBus_bits_data_6_1(WriteDataBuf_io_outputBus_bits_data_6_1),
    .io_outputBus_bits_data_6_2(WriteDataBuf_io_outputBus_bits_data_6_2),
    .io_outputBus_bits_data_6_3(WriteDataBuf_io_outputBus_bits_data_6_3),
    .io_outputBus_bits_data_7_0(WriteDataBuf_io_outputBus_bits_data_7_0),
    .io_outputBus_bits_data_7_1(WriteDataBuf_io_outputBus_bits_data_7_1),
    .io_outputBus_bits_data_7_2(WriteDataBuf_io_outputBus_bits_data_7_2),
    .io_outputBus_bits_data_7_3(WriteDataBuf_io_outputBus_bits_data_7_3),
    .io_outputBus_bits_instrId(WriteDataBuf_io_outputBus_bits_instrId),
    .io_wdbAlmostFull(WriteDataBuf_io_wdbAlmostFull)
  );
  Queue_50 coreRsp_Q ( // @[DCache.scala 96:25]
    .clock(coreRsp_Q_clock),
    .reset(coreRsp_Q_reset),
    .io_enq_ready(coreRsp_Q_io_enq_ready),
    .io_enq_valid(coreRsp_Q_io_enq_valid),
    .io_enq_bits_instrId(coreRsp_Q_io_enq_bits_instrId),
    .io_enq_bits_data_0(coreRsp_Q_io_enq_bits_data_0),
    .io_enq_bits_data_1(coreRsp_Q_io_enq_bits_data_1),
    .io_enq_bits_data_2(coreRsp_Q_io_enq_bits_data_2),
    .io_enq_bits_data_3(coreRsp_Q_io_enq_bits_data_3),
    .io_enq_bits_data_4(coreRsp_Q_io_enq_bits_data_4),
    .io_enq_bits_data_5(coreRsp_Q_io_enq_bits_data_5),
    .io_enq_bits_data_6(coreRsp_Q_io_enq_bits_data_6),
    .io_enq_bits_data_7(coreRsp_Q_io_enq_bits_data_7),
    .io_enq_bits_activeMask_0(coreRsp_Q_io_enq_bits_activeMask_0),
    .io_enq_bits_activeMask_1(coreRsp_Q_io_enq_bits_activeMask_1),
    .io_enq_bits_activeMask_2(coreRsp_Q_io_enq_bits_activeMask_2),
    .io_enq_bits_activeMask_3(coreRsp_Q_io_enq_bits_activeMask_3),
    .io_enq_bits_activeMask_4(coreRsp_Q_io_enq_bits_activeMask_4),
    .io_enq_bits_activeMask_5(coreRsp_Q_io_enq_bits_activeMask_5),
    .io_enq_bits_activeMask_6(coreRsp_Q_io_enq_bits_activeMask_6),
    .io_enq_bits_activeMask_7(coreRsp_Q_io_enq_bits_activeMask_7),
    .io_deq_ready(coreRsp_Q_io_deq_ready),
    .io_deq_valid(coreRsp_Q_io_deq_valid),
    .io_deq_bits_instrId(coreRsp_Q_io_deq_bits_instrId),
    .io_deq_bits_data_0(coreRsp_Q_io_deq_bits_data_0),
    .io_deq_bits_data_1(coreRsp_Q_io_deq_bits_data_1),
    .io_deq_bits_data_2(coreRsp_Q_io_deq_bits_data_2),
    .io_deq_bits_data_3(coreRsp_Q_io_deq_bits_data_3),
    .io_deq_bits_data_4(coreRsp_Q_io_deq_bits_data_4),
    .io_deq_bits_data_5(coreRsp_Q_io_deq_bits_data_5),
    .io_deq_bits_data_6(coreRsp_Q_io_deq_bits_data_6),
    .io_deq_bits_data_7(coreRsp_Q_io_deq_bits_data_7),
    .io_deq_bits_activeMask_0(coreRsp_Q_io_deq_bits_activeMask_0),
    .io_deq_bits_activeMask_1(coreRsp_Q_io_deq_bits_activeMask_1),
    .io_deq_bits_activeMask_2(coreRsp_Q_io_deq_bits_activeMask_2),
    .io_deq_bits_activeMask_3(coreRsp_Q_io_deq_bits_activeMask_3),
    .io_deq_bits_activeMask_4(coreRsp_Q_io_deq_bits_activeMask_4),
    .io_deq_bits_activeMask_5(coreRsp_Q_io_deq_bits_activeMask_5),
    .io_deq_bits_activeMask_6(coreRsp_Q_io_deq_bits_activeMask_6),
    .io_deq_bits_activeMask_7(coreRsp_Q_io_deq_bits_activeMask_7),
    .io_count(coreRsp_Q_io_count)
  );
  Queue_49 memRsp_Q ( // @[DCache.scala 99:24]
    .clock(memRsp_Q_clock),
    .reset(memRsp_Q_reset),
    .io_enq_ready(memRsp_Q_io_enq_ready),
    .io_enq_valid(memRsp_Q_io_enq_valid),
    .io_enq_bits_d_addr(memRsp_Q_io_enq_bits_d_addr),
    .io_enq_bits_d_data_0(memRsp_Q_io_enq_bits_d_data_0),
    .io_enq_bits_d_data_1(memRsp_Q_io_enq_bits_d_data_1),
    .io_enq_bits_d_data_2(memRsp_Q_io_enq_bits_d_data_2),
    .io_enq_bits_d_data_3(memRsp_Q_io_enq_bits_d_data_3),
    .io_enq_bits_d_data_4(memRsp_Q_io_enq_bits_d_data_4),
    .io_enq_bits_d_data_5(memRsp_Q_io_enq_bits_d_data_5),
    .io_enq_bits_d_data_6(memRsp_Q_io_enq_bits_d_data_6),
    .io_enq_bits_d_data_7(memRsp_Q_io_enq_bits_d_data_7),
    .io_deq_ready(memRsp_Q_io_deq_ready),
    .io_deq_valid(memRsp_Q_io_deq_valid),
    .io_deq_bits_d_addr(memRsp_Q_io_deq_bits_d_addr),
    .io_deq_bits_d_data_0(memRsp_Q_io_deq_bits_d_data_0),
    .io_deq_bits_d_data_1(memRsp_Q_io_deq_bits_d_data_1),
    .io_deq_bits_d_data_2(memRsp_Q_io_deq_bits_d_data_2),
    .io_deq_bits_d_data_3(memRsp_Q_io_deq_bits_d_data_3),
    .io_deq_bits_d_data_4(memRsp_Q_io_deq_bits_d_data_4),
    .io_deq_bits_d_data_5(memRsp_Q_io_deq_bits_d_data_5),
    .io_deq_bits_d_data_6(memRsp_Q_io_deq_bits_d_data_6),
    .io_deq_bits_d_data_7(memRsp_Q_io_deq_bits_d_data_7)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_clock),
    .reset(DataAccessesRRsp_DataAccess_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_1 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_1_clock),
    .reset(DataAccessesRRsp_DataAccess_1_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_1_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_1_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_1_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_1_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_1_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_1_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_1_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_1_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_1_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_2 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_2_clock),
    .reset(DataAccessesRRsp_DataAccess_2_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_2_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_2_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_2_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_2_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_2_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_2_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_2_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_2_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_2_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_3 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_3_clock),
    .reset(DataAccessesRRsp_DataAccess_3_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_3_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_3_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_3_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_3_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_3_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_3_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_3_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_3_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_3_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_4 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_4_clock),
    .reset(DataAccessesRRsp_DataAccess_4_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_4_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_4_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_4_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_4_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_4_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_4_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_4_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_4_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_4_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_5 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_5_clock),
    .reset(DataAccessesRRsp_DataAccess_5_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_5_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_5_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_5_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_5_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_5_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_5_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_5_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_5_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_5_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_6 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_6_clock),
    .reset(DataAccessesRRsp_DataAccess_6_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_6_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_6_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_6_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_6_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_6_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_6_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_6_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_6_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_6_io_w_req_bits_waymask)
  );
  SRAMTemplate_3 DataAccessesRRsp_DataAccess_7 ( // @[DCache.scala 240:28]
    .clock(DataAccessesRRsp_DataAccess_7_clock),
    .reset(DataAccessesRRsp_DataAccess_7_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_7_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_7_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_7_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_7_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_7_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_7_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_7_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_7_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_7_io_w_req_bits_waymask)
  );
  Arbiter_15 MemReqArb ( // @[DCache.scala 381:25]
    .io_in_0_ready(MemReqArb_io_in_0_ready),
    .io_in_0_valid(MemReqArb_io_in_0_valid),
    .io_in_0_bits_a_source(MemReqArb_io_in_0_bits_a_source),
    .io_in_0_bits_a_addr(MemReqArb_io_in_0_bits_a_addr),
    .io_in_1_ready(MemReqArb_io_in_1_ready),
    .io_in_1_valid(MemReqArb_io_in_1_valid),
    .io_in_1_bits_a_opcode(MemReqArb_io_in_1_bits_a_opcode),
    .io_in_1_bits_a_source(MemReqArb_io_in_1_bits_a_source),
    .io_in_1_bits_a_addr(MemReqArb_io_in_1_bits_a_addr),
    .io_in_1_bits_a_data_0(MemReqArb_io_in_1_bits_a_data_0),
    .io_in_1_bits_a_data_1(MemReqArb_io_in_1_bits_a_data_1),
    .io_in_1_bits_a_data_2(MemReqArb_io_in_1_bits_a_data_2),
    .io_in_1_bits_a_data_3(MemReqArb_io_in_1_bits_a_data_3),
    .io_in_1_bits_a_data_4(MemReqArb_io_in_1_bits_a_data_4),
    .io_in_1_bits_a_data_5(MemReqArb_io_in_1_bits_a_data_5),
    .io_in_1_bits_a_data_6(MemReqArb_io_in_1_bits_a_data_6),
    .io_in_1_bits_a_data_7(MemReqArb_io_in_1_bits_a_data_7),
    .io_in_1_bits_a_mask_0(MemReqArb_io_in_1_bits_a_mask_0),
    .io_in_1_bits_a_mask_1(MemReqArb_io_in_1_bits_a_mask_1),
    .io_in_1_bits_a_mask_2(MemReqArb_io_in_1_bits_a_mask_2),
    .io_in_1_bits_a_mask_3(MemReqArb_io_in_1_bits_a_mask_3),
    .io_in_1_bits_a_mask_4(MemReqArb_io_in_1_bits_a_mask_4),
    .io_in_1_bits_a_mask_5(MemReqArb_io_in_1_bits_a_mask_5),
    .io_in_1_bits_a_mask_6(MemReqArb_io_in_1_bits_a_mask_6),
    .io_in_1_bits_a_mask_7(MemReqArb_io_in_1_bits_a_mask_7),
    .io_out_ready(MemReqArb_io_out_ready),
    .io_out_valid(MemReqArb_io_out_valid),
    .io_out_bits_a_opcode(MemReqArb_io_out_bits_a_opcode),
    .io_out_bits_a_source(MemReqArb_io_out_bits_a_source),
    .io_out_bits_a_addr(MemReqArb_io_out_bits_a_addr),
    .io_out_bits_a_data_0(MemReqArb_io_out_bits_a_data_0),
    .io_out_bits_a_data_1(MemReqArb_io_out_bits_a_data_1),
    .io_out_bits_a_data_2(MemReqArb_io_out_bits_a_data_2),
    .io_out_bits_a_data_3(MemReqArb_io_out_bits_a_data_3),
    .io_out_bits_a_data_4(MemReqArb_io_out_bits_a_data_4),
    .io_out_bits_a_data_5(MemReqArb_io_out_bits_a_data_5),
    .io_out_bits_a_data_6(MemReqArb_io_out_bits_a_data_6),
    .io_out_bits_a_data_7(MemReqArb_io_out_bits_a_data_7),
    .io_out_bits_a_mask_0(MemReqArb_io_out_bits_a_mask_0),
    .io_out_bits_a_mask_1(MemReqArb_io_out_bits_a_mask_1),
    .io_out_bits_a_mask_2(MemReqArb_io_out_bits_a_mask_2),
    .io_out_bits_a_mask_3(MemReqArb_io_out_bits_a_mask_3),
    .io_out_bits_a_mask_4(MemReqArb_io_out_bits_a_mask_4),
    .io_out_bits_a_mask_5(MemReqArb_io_out_bits_a_mask_5),
    .io_out_bits_a_mask_6(MemReqArb_io_out_bits_a_mask_6),
    .io_out_bits_a_mask_7(MemReqArb_io_out_bits_a_mask_7)
  );
  assign io_coreReq_ready = _io_coreReq_ready_T_14 & MshrAccess_io_missReq_ready; // @[DCache.scala 340:42]
  assign io_coreRsp_valid = coreRsp_Q_io_deq_valid; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_instrId = coreRsp_Q_io_deq_bits_instrId; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_0 = coreRsp_Q_io_deq_bits_data_0; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_1 = coreRsp_Q_io_deq_bits_data_1; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_2 = coreRsp_Q_io_deq_bits_data_2; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_3 = coreRsp_Q_io_deq_bits_data_3; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_4 = coreRsp_Q_io_deq_bits_data_4; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_5 = coreRsp_Q_io_deq_bits_data_5; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_6 = coreRsp_Q_io_deq_bits_data_6; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_data_7 = coreRsp_Q_io_deq_bits_data_7; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_0 = coreRsp_Q_io_deq_bits_activeMask_0; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_1 = coreRsp_Q_io_deq_bits_activeMask_1; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_2 = coreRsp_Q_io_deq_bits_activeMask_2; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_3 = coreRsp_Q_io_deq_bits_activeMask_3; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_4 = coreRsp_Q_io_deq_bits_activeMask_4; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_5 = coreRsp_Q_io_deq_bits_activeMask_5; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_6 = coreRsp_Q_io_deq_bits_activeMask_6; // @[DCache.scala 314:20]
  assign io_coreRsp_bits_activeMask_7 = coreRsp_Q_io_deq_bits_activeMask_7; // @[DCache.scala 314:20]
  assign io_memRsp_ready = memRsp_Q_io_enq_ready; // @[DCache.scala 179:19]
  assign io_memReq_valid = MemReqArb_io_out_valid; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_opcode = MemReqArb_io_out_bits_a_opcode; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_source = MemReqArb_io_out_bits_a_source; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_addr = MemReqArb_io_out_bits_a_addr; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_0 = MemReqArb_io_out_bits_a_data_0; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_1 = MemReqArb_io_out_bits_a_data_1; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_2 = MemReqArb_io_out_bits_a_data_2; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_3 = MemReqArb_io_out_bits_a_data_3; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_4 = MemReqArb_io_out_bits_a_data_4; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_5 = MemReqArb_io_out_bits_a_data_5; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_6 = MemReqArb_io_out_bits_a_data_6; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_data_7 = MemReqArb_io_out_bits_a_data_7; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_0 = MemReqArb_io_out_bits_a_mask_0; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_1 = MemReqArb_io_out_bits_a_mask_1; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_2 = MemReqArb_io_out_bits_a_mask_2; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_3 = MemReqArb_io_out_bits_a_mask_3; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_4 = MemReqArb_io_out_bits_a_mask_4; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_5 = MemReqArb_io_out_bits_a_mask_5; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_6 = MemReqArb_io_out_bits_a_mask_6; // @[DCache.scala 402:13]
  assign io_memReq_bits_a_mask_7 = MemReqArb_io_out_bits_a_mask_7; // @[DCache.scala 402:13]
  assign BankConfArb_clock = clock;
  assign BankConfArb_reset = reset;
  assign BankConfArb_io_coreReqArb_isWrite = missRspFromMshr_st1 ? missRspTI_st1_isWrite : coreReq_st1_isWrite; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_enable = missRspFromMshr_st1 ? missRspFromMshr_st1 : cacheHit_st1; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_0_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_0_activeMask : coreReq_st1_perLaneAddr_0_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_0_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_0_blockOffset : coreReq_st1_perLaneAddr_0_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_0_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_0_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_1_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_1_activeMask : coreReq_st1_perLaneAddr_1_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_1_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_1_blockOffset : coreReq_st1_perLaneAddr_1_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_1_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_1_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_2_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_2_activeMask : coreReq_st1_perLaneAddr_2_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_2_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_2_blockOffset : coreReq_st1_perLaneAddr_2_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_2_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_2_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_3_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_3_activeMask : coreReq_st1_perLaneAddr_3_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_3_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_3_blockOffset : coreReq_st1_perLaneAddr_3_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_3_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_3_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_4_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_4_activeMask : coreReq_st1_perLaneAddr_4_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_4_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_4_blockOffset : coreReq_st1_perLaneAddr_4_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_4_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_4_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_5_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_5_activeMask : coreReq_st1_perLaneAddr_5_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_5_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_5_blockOffset : coreReq_st1_perLaneAddr_5_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_5_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_5_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_6_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_6_activeMask : coreReq_st1_perLaneAddr_6_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_6_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_6_blockOffset : coreReq_st1_perLaneAddr_6_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_6_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_6_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_7_activeMask = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_7_activeMask : coreReq_st1_perLaneAddr_7_activeMask; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_7_blockOffset = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_7_blockOffset : coreReq_st1_perLaneAddr_7_blockOffset; // @[DCache.scala 121:30]
  assign BankConfArb_io_coreReqArb_perLaneAddr_7_wordOffset1H = missRspFromMshr_st1 ?
    missRspTI_st1_perLaneAddr_7_wordOffset1H : 4'hf; // @[DCache.scala 121:30]
  assign MshrAccess_clock = clock;
  assign MshrAccess_reset = reset;
  assign MshrAccess_io_missReq_valid = cacheMiss_st1 & _MshrAccess_io_missReq_valid_T_2; // @[DCache.scala 191:48]
  assign MshrAccess_io_missReq_bits_blockAddr = {coreReq_st1_tag,coreReq_st1_setIdx}; // @[Cat.scala 31:58]
  assign MshrAccess_io_missReq_bits_instrId = coreReq_st1_instrId; // @[DCache.scala 197:38]
  assign MshrAccess_io_missReq_bits_targetInfo = {MshrAccess_io_missReq_bits_targetInfo_hi,
    MshrAccess_io_missReq_bits_targetInfo_lo}; // @[DCache.scala 199:64]
  assign MshrAccess_io_missRspIn_valid = memRsp_Q_io_deq_valid & _memRsp_Q_io_deq_ready_T_1; // @[DCache.scala 201:58]
  assign MshrAccess_io_missRspIn_bits_blockAddr = memRsp_Q_io_deq_bits_d_addr[31:5]; // @[L1CacheParameters.scala 55:41]
  assign MshrAccess_io_missRspOut_ready = _MshrAccess_io_missRspOut_ready_T_4 | _MshrAccess_io_missRspOut_ready_T_7; // @[DCache.scala 214:67]
  assign MshrAccess_io_miss2mem_ready = MemReqArb_io_in_0_ready; // @[DCache.scala 390:32]
  assign TagAccess_clock = clock;
  assign TagAccess_reset = reset;
  assign TagAccess_io_r_req_valid = io_coreReq_ready & io_coreReq_valid; // @[Decoupled.scala 50:35]
  assign TagAccess_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[DCache.scala 128:34]
  assign TagAccess_io_tagFromCore_st1 = coreReq_st1_tag; // @[DCache.scala 129:32]
  assign TagAccess_io_coreReqReady = io_coreReq_ready; // @[DCache.scala 130:29]
  assign TagAccess_io_w_req_valid = _missRspWriteEnable_T_3 & missRspFromMshr_st1 | _T_5; // @[DCache.scala 233:73]
  assign TagAccess_io_w_req_bits_setIdx = memRsp_Q_io_deq_bits_d_addr[9:5]; // @[L1CacheParameters.scala 45:9]
  assign TagAccess_io_w_req_bits_data_0 = memRsp_Q_io_deq_bits_d_addr[31:10]; // @[L1CacheParameters.scala 43:35]
  assign TagAccess_io_w_req_bits_data_1 = memRsp_Q_io_deq_bits_d_addr[31:10]; // @[L1CacheParameters.scala 43:35]
  assign DataCorssBar_io_DataIn_0 = readMissRsp_st2 ? r_0_0 : _T_14_0; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_1 = readMissRsp_st2 ? r_0_1 : _T_14_1; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_2 = readMissRsp_st2 ? r_0_2 : _T_14_2; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_3 = readMissRsp_st2 ? r_0_3 : _T_14_3; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_4 = readMissRsp_st2 ? r_0_4 : _T_14_4; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_5 = readMissRsp_st2 ? r_0_5 : _T_14_5; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_6 = readMissRsp_st2 ? r_0_6 : _T_14_6; // @[DCache.scala 301:32]
  assign DataCorssBar_io_DataIn_7 = readMissRsp_st2 ? r_0_7 : _T_14_7; // @[DCache.scala 301:32]
  assign DataCorssBar_io_Select1H_0 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_0 :
    arbDataCrsbarSel1H_st3_0; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_1 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_1 :
    arbDataCrsbarSel1H_st3_1; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_2 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_2 :
    arbDataCrsbarSel1H_st3_2; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_3 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_3 :
    arbDataCrsbarSel1H_st3_3; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_4 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_4 :
    arbDataCrsbarSel1H_st3_4; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_5 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_5 :
    arbDataCrsbarSel1H_st3_5; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_6 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_6 :
    arbDataCrsbarSel1H_st3_6; // @[DCache.scala 308:34]
  assign DataCorssBar_io_Select1H_7 = coreReq_st2_isWrite | readMissRsp_st2 ? arbDataCrsbarSel1H_st2_7 :
    arbDataCrsbarSel1H_st3_7; // @[DCache.scala 308:34]
  assign WriteDataBuf_clock = clock;
  assign WriteDataBuf_reset = reset;
  assign WriteDataBuf_io_inputBus_valid = writeMiss_st2 | writeHit_st2 | _WriteDataBuf_io_inputBus_valid_T_1; // @[DCache.scala 344:66]
  assign WriteDataBuf_io_inputBus_bits_mask_0 = arbArrayEn_st2_0 ? _WriteDataBuf_io_inputBus_bits_mask_0_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_1 = arbArrayEn_st2_1 ? _WriteDataBuf_io_inputBus_bits_mask_1_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_2 = arbArrayEn_st2_2 ? _WriteDataBuf_io_inputBus_bits_mask_2_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_3 = arbArrayEn_st2_3 ? _WriteDataBuf_io_inputBus_bits_mask_3_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_4 = arbArrayEn_st2_4 ? _WriteDataBuf_io_inputBus_bits_mask_4_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_5 = arbArrayEn_st2_5 ? _WriteDataBuf_io_inputBus_bits_mask_5_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_6 = arbArrayEn_st2_6 ? _WriteDataBuf_io_inputBus_bits_mask_6_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_mask_7 = arbArrayEn_st2_7 ? _WriteDataBuf_io_inputBus_bits_mask_7_T_2 : 4'h0; // @[DCache.scala 358:12]
  assign WriteDataBuf_io_inputBus_bits_addr = {WriteDataBuf_io_inputBus_bits_addr_hi,5'h0}; // @[Cat.scala 31:58]
  assign WriteDataBuf_io_inputBus_bits_data_0_0 = arbArrayEn_st2_0 ? _WriteDataBuf_io_inputBus_bits_data_0_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_0_1 = arbArrayEn_st2_0 ? _WriteDataBuf_io_inputBus_bits_data_0_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_0_2 = arbArrayEn_st2_0 ? _WriteDataBuf_io_inputBus_bits_data_0_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_0_3 = arbArrayEn_st2_0 ? _WriteDataBuf_io_inputBus_bits_data_0_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_1_0 = arbArrayEn_st2_1 ? _WriteDataBuf_io_inputBus_bits_data_1_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_1_1 = arbArrayEn_st2_1 ? _WriteDataBuf_io_inputBus_bits_data_1_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_1_2 = arbArrayEn_st2_1 ? _WriteDataBuf_io_inputBus_bits_data_1_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_1_3 = arbArrayEn_st2_1 ? _WriteDataBuf_io_inputBus_bits_data_1_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_2_0 = arbArrayEn_st2_2 ? _WriteDataBuf_io_inputBus_bits_data_2_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_2_1 = arbArrayEn_st2_2 ? _WriteDataBuf_io_inputBus_bits_data_2_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_2_2 = arbArrayEn_st2_2 ? _WriteDataBuf_io_inputBus_bits_data_2_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_2_3 = arbArrayEn_st2_2 ? _WriteDataBuf_io_inputBus_bits_data_2_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_3_0 = arbArrayEn_st2_3 ? _WriteDataBuf_io_inputBus_bits_data_3_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_3_1 = arbArrayEn_st2_3 ? _WriteDataBuf_io_inputBus_bits_data_3_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_3_2 = arbArrayEn_st2_3 ? _WriteDataBuf_io_inputBus_bits_data_3_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_3_3 = arbArrayEn_st2_3 ? _WriteDataBuf_io_inputBus_bits_data_3_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_4_0 = arbArrayEn_st2_4 ? _WriteDataBuf_io_inputBus_bits_data_4_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_4_1 = arbArrayEn_st2_4 ? _WriteDataBuf_io_inputBus_bits_data_4_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_4_2 = arbArrayEn_st2_4 ? _WriteDataBuf_io_inputBus_bits_data_4_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_4_3 = arbArrayEn_st2_4 ? _WriteDataBuf_io_inputBus_bits_data_4_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_5_0 = arbArrayEn_st2_5 ? _WriteDataBuf_io_inputBus_bits_data_5_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_5_1 = arbArrayEn_st2_5 ? _WriteDataBuf_io_inputBus_bits_data_5_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_5_2 = arbArrayEn_st2_5 ? _WriteDataBuf_io_inputBus_bits_data_5_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_5_3 = arbArrayEn_st2_5 ? _WriteDataBuf_io_inputBus_bits_data_5_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_6_0 = arbArrayEn_st2_6 ? _WriteDataBuf_io_inputBus_bits_data_6_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_6_1 = arbArrayEn_st2_6 ? _WriteDataBuf_io_inputBus_bits_data_6_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_6_2 = arbArrayEn_st2_6 ? _WriteDataBuf_io_inputBus_bits_data_6_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_6_3 = arbArrayEn_st2_6 ? _WriteDataBuf_io_inputBus_bits_data_6_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_7_0 = arbArrayEn_st2_7 ? _WriteDataBuf_io_inputBus_bits_data_7_0_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_7_1 = arbArrayEn_st2_7 ? _WriteDataBuf_io_inputBus_bits_data_7_1_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_7_2 = arbArrayEn_st2_7 ? _WriteDataBuf_io_inputBus_bits_data_7_2_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_data_7_3 = arbArrayEn_st2_7 ? _WriteDataBuf_io_inputBus_bits_data_7_3_T_3 : 8'h0; // @[DCache.scala 365:14]
  assign WriteDataBuf_io_inputBus_bits_instrId = coreReq_st2_instrId; // @[DCache.scala 374:41]
  assign WriteDataBuf_io_inputBus_bits_bankConflict = bankConflict_st2; // @[DCache.scala 376:46]
  assign WriteDataBuf_io_inputBus_bits_subWordMissReq = writeMissSubWord_st2; // @[DCache.scala 377:48]
  assign WriteDataBuf_io_inputBus_bits_subWordMissRsp = writeMissRsp_st2 & missRspTI_st1_isWrite; // @[DCache.scala 378:68]
  assign WriteDataBuf_io_outputBus_ready = MemReqArb_io_in_1_ready; // @[DCache.scala 399:35]
  assign coreRsp_Q_clock = clock;
  assign coreRsp_Q_reset = reset;
  assign coreRsp_Q_io_enq_valid = readHit_st3 | readMissRsp_st2 | writeMiss_st3 | writeHit_st3; // @[DCache.scala 315:77]
  assign coreRsp_Q_io_enq_bits_instrId = readMissRsp_st2 ? memRspInstrId_st2 : coreReqInstrId_st3; // @[DCache.scala 322:39]
  assign coreRsp_Q_io_enq_bits_data_0 = DataCorssBar_io_DataOut_0; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_1 = DataCorssBar_io_DataOut_1; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_2 = DataCorssBar_io_DataOut_2; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_3 = DataCorssBar_io_DataOut_3; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_4 = DataCorssBar_io_DataOut_4; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_5 = DataCorssBar_io_DataOut_5; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_6 = DataCorssBar_io_DataOut_6; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_data_7 = DataCorssBar_io_DataOut_7; // @[DCache.scala 321:30]
  assign coreRsp_Q_io_enq_bits_activeMask_0 = readMissRsp_st2 ? missRspTILaneMask_st2_0 : coreReqActvMask_st3_0; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_1 = readMissRsp_st2 ? missRspTILaneMask_st2_1 : coreReqActvMask_st3_1; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_2 = readMissRsp_st2 ? missRspTILaneMask_st2_2 : coreReqActvMask_st3_2; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_3 = readMissRsp_st2 ? missRspTILaneMask_st2_3 : coreReqActvMask_st3_3; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_4 = readMissRsp_st2 ? missRspTILaneMask_st2_4 : coreReqActvMask_st3_4; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_5 = readMissRsp_st2 ? missRspTILaneMask_st2_5 : coreReqActvMask_st3_5; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_6 = readMissRsp_st2 ? missRspTILaneMask_st2_6 : coreReqActvMask_st3_6; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_enq_bits_activeMask_7 = readMissRsp_st2 ? missRspTILaneMask_st2_7 : coreReqActvMask_st3_7; // @[DCache.scala 327:42]
  assign coreRsp_Q_io_deq_ready = io_coreRsp_ready; // @[DCache.scala 314:20]
  assign memRsp_Q_clock = clock;
  assign memRsp_Q_reset = reset;
  assign memRsp_Q_io_enq_valid = io_memRsp_valid; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_addr = io_memRsp_bits_d_addr; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_0 = io_memRsp_bits_d_data_0; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_1 = io_memRsp_bits_d_data_1; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_2 = io_memRsp_bits_d_data_2; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_3 = io_memRsp_bits_d_data_3; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_4 = io_memRsp_bits_d_data_4; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_5 = io_memRsp_bits_d_data_5; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_6 = io_memRsp_bits_d_data_6; // @[DCache.scala 179:19]
  assign memRsp_Q_io_enq_bits_d_data_7 = io_memRsp_bits_d_data_7; // @[DCache.scala 179:19]
  assign memRsp_Q_io_deq_ready = MshrAccess_io_missRspIn_ready & ~(readHit_st2 | writeHit_st2); // @[DCache.scala 180:58]
  assign DataAccessesRRsp_DataAccess_clock = clock;
  assign DataAccessesRRsp_DataAccess_reset = reset;
  assign DataAccessesRRsp_DataAccess_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_0 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_2; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_io_w_req_valid = missRspWriteEnable | _DataAccessesRRsp_DataAccess_io_w_req_valid_T
    ; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_0 = _DataAccessesRRsp_T__0[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_1 = _DataAccessesRRsp_T__0[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_2 = _DataAccessesRRsp_T__0[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_3 = _DataAccessesRRsp_T__0[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_0_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_1_clock = clock;
  assign DataAccessesRRsp_DataAccess_1_reset = reset;
  assign DataAccessesRRsp_DataAccess_1_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_1 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_6; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_1_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_2; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_0 = _DataAccessesRRsp_T__1[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_1 = _DataAccessesRRsp_T__1[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_2 = _DataAccessesRRsp_T__1[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_3 = _DataAccessesRRsp_T__1[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_1_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_2_clock = clock;
  assign DataAccessesRRsp_DataAccess_2_reset = reset;
  assign DataAccessesRRsp_DataAccess_2_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_2 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_10; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_2_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_4; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_0 = _DataAccessesRRsp_T__2[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_1 = _DataAccessesRRsp_T__2[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_2 = _DataAccessesRRsp_T__2[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_3 = _DataAccessesRRsp_T__2[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_2_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_3_clock = clock;
  assign DataAccessesRRsp_DataAccess_3_reset = reset;
  assign DataAccessesRRsp_DataAccess_3_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_3 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_14; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_3_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_6; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_0 = _DataAccessesRRsp_T__3[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_1 = _DataAccessesRRsp_T__3[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_2 = _DataAccessesRRsp_T__3[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_3 = _DataAccessesRRsp_T__3[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_3_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_4_clock = clock;
  assign DataAccessesRRsp_DataAccess_4_reset = reset;
  assign DataAccessesRRsp_DataAccess_4_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_4 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_18; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_4_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_8; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_0 = _DataAccessesRRsp_T__4[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_1 = _DataAccessesRRsp_T__4[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_2 = _DataAccessesRRsp_T__4[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_3 = _DataAccessesRRsp_T__4[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_4_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_5_clock = clock;
  assign DataAccessesRRsp_DataAccess_5_reset = reset;
  assign DataAccessesRRsp_DataAccess_5_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_5 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_22; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_5_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_10; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_0 = _DataAccessesRRsp_T__5[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_1 = _DataAccessesRRsp_T__5[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_2 = _DataAccessesRRsp_T__5[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_3 = _DataAccessesRRsp_T__5[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_5_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_6_clock = clock;
  assign DataAccessesRRsp_DataAccess_6_reset = reset;
  assign DataAccessesRRsp_DataAccess_6_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_6 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_26; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_6_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_12; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_0 = _DataAccessesRRsp_T__6[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_1 = _DataAccessesRRsp_T__6[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_2 = _DataAccessesRRsp_T__6[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_3 = _DataAccessesRRsp_T__6[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_6_wordOffset1H; // @[DCache.scala 279:54]
  assign DataAccessesRRsp_DataAccess_7_clock = clock;
  assign DataAccessesRRsp_DataAccess_7_reset = reset;
  assign DataAccessesRRsp_DataAccess_7_io_r_req_valid = readHit_st1 & BankConfArb_io_dataArrayEn_7 |
    _DataAccessesRRsp_DataAccess_io_r_req_valid_T_30; // @[DCache.scala 285:80]
  assign DataAccessesRRsp_DataAccess_7_io_r_req_bits_setIdx = {coreReq_st1_setIdx,wayIdxAtHit_st1}; // @[Cat.scala 31:58]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_valid = missRspWriteEnable |
    _DataAccessesRRsp_DataAccess_io_w_req_valid_T_14; // @[DCache.scala 248:37]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_setIdx = missRspWriteEnable ?
    DataAccessesRRsp_DAWtSetIdxMissRspCase_st1 : DataAccessesRRsp_DAWtSetIdxWtHitCase_st2; // @[DCache.scala 274:43]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_0 = _DataAccessesRRsp_T__7[7:0]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_1 = _DataAccessesRRsp_T__7[15:8]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_2 = _DataAccessesRRsp_T__7[23:16]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_3 = _DataAccessesRRsp_T__7[31:24]; // @[DCache.scala 256:73]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_waymask = missRspWriteEnable ? 4'hf :
    arbAddrCrsbarOut_st2_7_wordOffset1H; // @[DCache.scala 279:54]
  assign MemReqArb_io_in_0_valid = MshrAccess_io_miss2mem_valid; // @[DCache.scala 403:28]
  assign MemReqArb_io_in_0_bits_a_source = MshrAccess_io_miss2mem_bits_instrId; // @[DCache.scala 384:24 388:23]
  assign MemReqArb_io_in_0_bits_a_addr = {MshrAccess_io_miss2mem_bits_blockAddr,5'h0}; // @[Cat.scala 31:58]
  assign MemReqArb_io_in_1_valid = WriteDataBuf_io_outputBus_valid; // @[DCache.scala 405:28]
  assign MemReqArb_io_in_1_bits_a_opcode = &_wdbMemReq_a_opcode_T ? 3'h0 : 3'h1; // @[DCache.scala 394:28]
  assign MemReqArb_io_in_1_bits_a_source = WriteDataBuf_io_outputBus_bits_instrId; // @[DCache.scala 392:23 397:22]
  assign MemReqArb_io_in_1_bits_a_addr = WriteDataBuf_io_outputBus_bits_addr; // @[DCache.scala 392:23 395:20]
  assign MemReqArb_io_in_1_bits_a_data_0 = _T_52[31:0]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_1 = _T_52[63:32]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_2 = _T_52[95:64]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_3 = _T_52[127:96]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_4 = _T_52[159:128]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_5 = _T_52[191:160]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_6 = _T_52[223:192]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_data_7 = _T_52[255:224]; // @[DCache.scala 396:48]
  assign MemReqArb_io_in_1_bits_a_mask_0 = WriteDataBuf_io_outputBus_bits_mask_0; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_1 = WriteDataBuf_io_outputBus_bits_mask_1; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_2 = WriteDataBuf_io_outputBus_bits_mask_2; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_3 = WriteDataBuf_io_outputBus_bits_mask_3; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_4 = WriteDataBuf_io_outputBus_bits_mask_4; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_5 = WriteDataBuf_io_outputBus_bits_mask_5; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_6 = WriteDataBuf_io_outputBus_bits_mask_6; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_in_1_bits_a_mask_7 = WriteDataBuf_io_outputBus_bits_mask_7; // @[DCache.scala 392:23 398:20]
  assign MemReqArb_io_out_ready = io_memReq_ready; // @[DCache.scala 402:13]
  always @(posedge clock) begin
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_instrId <= io_coreReq_bits_instrId; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_isWrite <= io_coreReq_bits_isWrite; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_tag <= io_coreReq_bits_tag; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_setIdx <= io_coreReq_bits_setIdx; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_0_activeMask <= io_coreReq_bits_perLaneAddr_0_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_0_blockOffset <= io_coreReq_bits_perLaneAddr_0_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_1_activeMask <= io_coreReq_bits_perLaneAddr_1_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_1_blockOffset <= io_coreReq_bits_perLaneAddr_1_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_2_activeMask <= io_coreReq_bits_perLaneAddr_2_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_2_blockOffset <= io_coreReq_bits_perLaneAddr_2_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_3_activeMask <= io_coreReq_bits_perLaneAddr_3_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_3_blockOffset <= io_coreReq_bits_perLaneAddr_3_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_4_activeMask <= io_coreReq_bits_perLaneAddr_4_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_4_blockOffset <= io_coreReq_bits_perLaneAddr_4_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_5_activeMask <= io_coreReq_bits_perLaneAddr_5_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_5_blockOffset <= io_coreReq_bits_perLaneAddr_5_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_6_activeMask <= io_coreReq_bits_perLaneAddr_6_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_6_blockOffset <= io_coreReq_bits_perLaneAddr_6_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_7_activeMask <= io_coreReq_bits_perLaneAddr_7_activeMask; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_7_blockOffset <= io_coreReq_bits_perLaneAddr_7_blockOffset; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_0 <= io_coreReq_bits_data_0; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_1 <= io_coreReq_bits_data_1; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_2 <= io_coreReq_bits_data_2; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_3 <= io_coreReq_bits_data_3; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_4 <= io_coreReq_bits_data_4; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_5 <= io_coreReq_bits_data_5; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_6 <= io_coreReq_bits_data_6; // @[Reg.scala 17:22]
    end
    if (_coreReq_st1_T) begin // @[Reg.scala 17:18]
      coreReq_st1_data_7 <= io_coreReq_bits_data_7; // @[Reg.scala 17:22]
    end
    coreReq_st2_instrId <= coreReq_st1_instrId; // @[DCache.scala 105:28]
    coreReq_st2_isWrite <= coreReq_st1_isWrite; // @[DCache.scala 105:28]
    coreReq_st2_tag <= coreReq_st1_tag; // @[DCache.scala 105:28]
    coreReq_st2_setIdx <= coreReq_st1_setIdx; // @[DCache.scala 105:28]
    coreReq_st2_data_0 <= coreReq_st1_data_0; // @[DCache.scala 105:28]
    coreReq_st2_data_1 <= coreReq_st1_data_1; // @[DCache.scala 105:28]
    coreReq_st2_data_2 <= coreReq_st1_data_2; // @[DCache.scala 105:28]
    coreReq_st2_data_3 <= coreReq_st1_data_3; // @[DCache.scala 105:28]
    coreReq_st2_data_4 <= coreReq_st1_data_4; // @[DCache.scala 105:28]
    coreReq_st2_data_5 <= coreReq_st1_data_5; // @[DCache.scala 105:28]
    coreReq_st2_data_6 <= coreReq_st1_data_6; // @[DCache.scala 105:28]
    coreReq_st2_data_7 <= coreReq_st1_data_7; // @[DCache.scala 105:28]
    coreReqInstrId_st3 <= coreReq_st2_instrId; // @[DCache.scala 106:35]
    coreReqActvMask_st3_r_0 <= BankConfArb_io_activeLane_0; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_1 <= BankConfArb_io_activeLane_1; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_2 <= BankConfArb_io_activeLane_2; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_3 <= BankConfArb_io_activeLane_3; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_4 <= BankConfArb_io_activeLane_4; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_5 <= BankConfArb_io_activeLane_5; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_6 <= BankConfArb_io_activeLane_6; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_r_7 <= BankConfArb_io_activeLane_7; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_0 <= coreReqActvMask_st3_r_0; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_1 <= coreReqActvMask_st3_r_1; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_2 <= coreReqActvMask_st3_r_2; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_3 <= coreReqActvMask_st3_r_3; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_4 <= coreReqActvMask_st3_r_4; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_5 <= coreReqActvMask_st3_r_5; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_6 <= coreReqActvMask_st3_r_6; // @[Reg.scala 16:16 17:{18,22}]
    coreReqActvMask_st3_7 <= coreReqActvMask_st3_r_7; // @[Reg.scala 16:16 17:{18,22}]
    cacheHit_st1_REG <= io_coreReq_ready & io_coreReq_valid; // @[Decoupled.scala 50:35]
    if (MshrAccess_io_missReq_ready) begin // @[Reg.scala 17:18]
      cacheMiss_st1_r <= _coreReq_st1_T; // @[Reg.scala 17:22]
    end
    wayIdxAtHit_st2 <= TagAccess_io_waymaskHit_st1[1]; // @[CircuitMath.scala 30:8]
    writeMiss_st2 <= cacheMiss_st1 & coreReq_st1_isWrite; // @[DCache.scala 156:37]
    writeMissSubWord_st2 <= writeMiss_st1 & byteEn_st1; // @[DCache.scala 158:44]
    writeMiss_st3 <= writeMiss_st2; // @[DCache.scala 162:30]
    if (reset) begin // @[DCache.scala 164:28]
      readHit_st2 <= 1'h0; // @[DCache.scala 164:28]
    end else begin
      readHit_st2 <= readHit_st1 | readHit_st2 & readHit_st2_REG; // @[DCache.scala 165:15]
    end
    readHit_st2_REG <= BankConfArb_io_bankConflict; // @[DCache.scala 165:56]
    readHit_st3 <= readHit_st2; // @[DCache.scala 167:28]
    writeHit_st2 <= cacheHit_st1 & coreReq_st1_isWrite; // @[DCache.scala 155:35]
    writeHit_st3 <= writeHit_st2; // @[DCache.scala 169:29]
    bankConflict_st2 <= BankConfArb_io_bankConflict; // @[DCache.scala 171:33]
    arbDataCrsbarSel1H_st2_0 <= BankConfArb_io_dataCrsbarSel1H_0; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_1 <= BankConfArb_io_dataCrsbarSel1H_1; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_2 <= BankConfArb_io_dataCrsbarSel1H_2; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_3 <= BankConfArb_io_dataCrsbarSel1H_3; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_4 <= BankConfArb_io_dataCrsbarSel1H_4; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_5 <= BankConfArb_io_dataCrsbarSel1H_5; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_6 <= BankConfArb_io_dataCrsbarSel1H_6; // @[DCache.scala 172:39]
    arbDataCrsbarSel1H_st2_7 <= BankConfArb_io_dataCrsbarSel1H_7; // @[DCache.scala 172:39]
    arbAddrCrsbarOut_st2_0_wordOffset1H <= BankConfArb_io_addrCrsbarOut_0_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_1_wordOffset1H <= BankConfArb_io_addrCrsbarOut_1_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_2_wordOffset1H <= BankConfArb_io_addrCrsbarOut_2_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_3_wordOffset1H <= BankConfArb_io_addrCrsbarOut_3_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_4_wordOffset1H <= BankConfArb_io_addrCrsbarOut_4_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_5_wordOffset1H <= BankConfArb_io_addrCrsbarOut_5_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_6_wordOffset1H <= BankConfArb_io_addrCrsbarOut_6_wordOffset1H; // @[DCache.scala 173:37]
    arbAddrCrsbarOut_st2_7_wordOffset1H <= BankConfArb_io_addrCrsbarOut_7_wordOffset1H; // @[DCache.scala 173:37]
    arbArrayEn_st2_0 <= BankConfArb_io_dataArrayEn_0; // @[DCache.scala 174:31]
    arbArrayEn_st2_1 <= BankConfArb_io_dataArrayEn_1; // @[DCache.scala 174:31]
    arbArrayEn_st2_2 <= BankConfArb_io_dataArrayEn_2; // @[DCache.scala 174:31]
    arbArrayEn_st2_3 <= BankConfArb_io_dataArrayEn_3; // @[DCache.scala 174:31]
    arbArrayEn_st2_4 <= BankConfArb_io_dataArrayEn_4; // @[DCache.scala 174:31]
    arbArrayEn_st2_5 <= BankConfArb_io_dataArrayEn_5; // @[DCache.scala 174:31]
    arbArrayEn_st2_6 <= BankConfArb_io_dataArrayEn_6; // @[DCache.scala 174:31]
    arbArrayEn_st2_7 <= BankConfArb_io_dataArrayEn_7; // @[DCache.scala 174:31]
    arbDataCrsbarSel1H_st3_0 <= arbDataCrsbarSel1H_st2_0; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_1 <= arbDataCrsbarSel1H_st2_1; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_2 <= arbDataCrsbarSel1H_st2_2; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_3 <= arbDataCrsbarSel1H_st2_3; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_4 <= arbDataCrsbarSel1H_st2_4; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_5 <= arbDataCrsbarSel1H_st2_5; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_6 <= arbDataCrsbarSel1H_st2_6; // @[DCache.scala 176:39]
    arbDataCrsbarSel1H_st3_7 <= arbDataCrsbarSel1H_st2_7; // @[DCache.scala 176:39]
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_0 <= memRspData_st1_0_0; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_1 <= memRspData_st1_0_1; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_2 <= memRspData_st1_0_2; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_3 <= memRspData_st1_0_3; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_4 <= memRspData_st1_0_4; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_5 <= memRspData_st1_0_5; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_6 <= memRspData_st1_0_6; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      r_0_7 <= memRspData_st1_0_7; // @[Reg.scala 17:22]
    end
    missRspTILaneMask_st2_0 <= BankConfArb_io_activeLane_0; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_1 <= BankConfArb_io_activeLane_1; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_2 <= BankConfArb_io_activeLane_2; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_3 <= BankConfArb_io_activeLane_3; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_4 <= BankConfArb_io_activeLane_4; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_5 <= BankConfArb_io_activeLane_5; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_6 <= BankConfArb_io_activeLane_6; // @[DCache.scala 207:38]
    missRspTILaneMask_st2_7 <= BankConfArb_io_activeLane_7; // @[DCache.scala 207:38]
    memRspInstrId_st2 <= MshrAccess_io_missRspOut_bits_instrId; // @[DCache.scala 208:34]
    if (_T_11) begin // @[DCache.scala 227:73]
      readMissRspCnter <= 1'h0; // @[DCache.scala 228:22]
    end else if (missRspFromMshr_st1 & _T_5) begin // @[DCache.scala 229:75]
      readMissRspCnter <= readMissRspCnter + 1'h1; // @[DCache.scala 230:22]
    end
    readMissRsp_st2 <= (_readMissRsp_st1_T | MshrAccess_io_missRspOut_valid & BankConfArb_io_bankConflict) &
      _MshrAccess_io_missRspOut_ready_T; // @[DCache.scala 220:126]
    writeMissRsp_st2 <= _readMissRsp_st1_T & missRspTI_st1_isWrite; // @[DCache.scala 221:58]
    REG <= MshrAccess_io_missRspOut_valid; // @[DCache.scala 204:23 88:33]
    REG_1 <= MshrAccess_io_missRspOut_bits_blockAddr; // @[DCache.scala 227:13]
    missRspWriteEnable_REG <= MshrAccess_io_missRspOut_valid; // @[DCache.scala 204:23 88:33]
    missRspWriteEnable_REG_1 <= MshrAccess_io_missRspOut_bits_blockAddr; // @[DCache.scala 233:13]
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_0 <= DataAccessesRRsp_0; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_1 <= DataAccessesRRsp_1; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_2 <= DataAccessesRRsp_2; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_3 <= DataAccessesRRsp_3; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_4 <= DataAccessesRRsp_4; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_5 <= DataAccessesRRsp_5; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_6 <= DataAccessesRRsp_6; // @[Reg.scala 17:22]
    end
    if (readHit_st2) begin // @[Reg.scala 17:18]
      dataAccess_data_st3_7 <= DataAccessesRRsp_7; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  coreReq_st1_instrId = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  coreReq_st1_isWrite = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  coreReq_st1_tag = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  coreReq_st1_setIdx = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_0_activeMask = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_0_blockOffset = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_1_activeMask = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_1_blockOffset = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_2_activeMask = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_2_blockOffset = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_3_activeMask = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_3_blockOffset = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_4_activeMask = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_4_blockOffset = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_5_activeMask = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_5_blockOffset = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_6_activeMask = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_6_blockOffset = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_7_activeMask = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_7_blockOffset = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  coreReq_st1_data_0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  coreReq_st1_data_1 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  coreReq_st1_data_2 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  coreReq_st1_data_3 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  coreReq_st1_data_4 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  coreReq_st1_data_5 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  coreReq_st1_data_6 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  coreReq_st1_data_7 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  coreReq_st2_instrId = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  coreReq_st2_isWrite = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  coreReq_st2_tag = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  coreReq_st2_setIdx = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  coreReq_st2_data_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  coreReq_st2_data_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  coreReq_st2_data_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  coreReq_st2_data_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  coreReq_st2_data_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  coreReq_st2_data_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  coreReq_st2_data_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  coreReq_st2_data_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  coreReqInstrId_st3 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  coreReqActvMask_st3_r_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  coreReqActvMask_st3_r_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  coreReqActvMask_st3_r_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  coreReqActvMask_st3_r_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  coreReqActvMask_st3_r_4 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  coreReqActvMask_st3_r_5 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  coreReqActvMask_st3_r_6 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  coreReqActvMask_st3_r_7 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  coreReqActvMask_st3_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  coreReqActvMask_st3_1 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  coreReqActvMask_st3_2 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  coreReqActvMask_st3_3 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  coreReqActvMask_st3_4 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  coreReqActvMask_st3_5 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  coreReqActvMask_st3_6 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  coreReqActvMask_st3_7 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  cacheHit_st1_REG = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  cacheMiss_st1_r = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  wayIdxAtHit_st2 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  writeMiss_st2 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  writeMissSubWord_st2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  writeMiss_st3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  readHit_st2 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  readHit_st2_REG = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  readHit_st3 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  writeHit_st2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  writeHit_st3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  bankConflict_st2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_0 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_1 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_2 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_3 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_4 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_5 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_6 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_7 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_0_wordOffset1H = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_1_wordOffset1H = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_2_wordOffset1H = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_3_wordOffset1H = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_4_wordOffset1H = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_5_wordOffset1H = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_6_wordOffset1H = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  arbAddrCrsbarOut_st2_7_wordOffset1H = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  arbArrayEn_st2_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  arbArrayEn_st2_1 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  arbArrayEn_st2_2 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  arbArrayEn_st2_3 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  arbArrayEn_st2_4 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  arbArrayEn_st2_5 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  arbArrayEn_st2_6 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  arbArrayEn_st2_7 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_0 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_1 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_2 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_3 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_4 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_5 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_6 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st3_7 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  r_0_0 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  r_0_1 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  r_0_2 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  r_0_3 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  r_0_4 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  r_0_5 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  r_0_6 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  r_0_7 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  missRspTILaneMask_st2_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  missRspTILaneMask_st2_1 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  missRspTILaneMask_st2_2 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  missRspTILaneMask_st2_3 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  missRspTILaneMask_st2_4 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  missRspTILaneMask_st2_5 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  missRspTILaneMask_st2_6 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  missRspTILaneMask_st2_7 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  memRspInstrId_st2 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  readMissRspCnter = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  readMissRsp_st2 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  writeMissRsp_st2 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  REG = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  REG_1 = _RAND_122[26:0];
  _RAND_123 = {1{`RANDOM}};
  missRspWriteEnable_REG = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  missRspWriteEnable_REG_1 = _RAND_124[26:0];
  _RAND_125 = {1{`RANDOM}};
  dataAccess_data_st3_0 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  dataAccess_data_st3_1 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  dataAccess_data_st3_2 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  dataAccess_data_st3_3 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  dataAccess_data_st3_4 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  dataAccess_data_st3_5 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  dataAccess_data_st3_6 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  dataAccess_data_st3_7 = _RAND_132[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BankConflictArbiter_1(
  input        clock,
  input        reset,
  input        io_coreReqArb_isWrite,
  input        io_coreReqArb_perLaneAddr_0_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_0_blockOffset,
  input        io_coreReqArb_perLaneAddr_1_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_1_blockOffset,
  input        io_coreReqArb_perLaneAddr_2_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_2_blockOffset,
  input        io_coreReqArb_perLaneAddr_3_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_3_blockOffset,
  input        io_coreReqArb_perLaneAddr_4_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_4_blockOffset,
  input        io_coreReqArb_perLaneAddr_5_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_5_blockOffset,
  input        io_coreReqArb_perLaneAddr_6_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_6_blockOffset,
  input        io_coreReqArb_perLaneAddr_7_activeMask,
  input  [2:0] io_coreReqArb_perLaneAddr_7_blockOffset,
  output [7:0] io_dataCrsbarSel1H_0,
  output [7:0] io_dataCrsbarSel1H_1,
  output [7:0] io_dataCrsbarSel1H_2,
  output [7:0] io_dataCrsbarSel1H_3,
  output [7:0] io_dataCrsbarSel1H_4,
  output [7:0] io_dataCrsbarSel1H_5,
  output [7:0] io_dataCrsbarSel1H_6,
  output [7:0] io_dataCrsbarSel1H_7,
  output [3:0] io_addrCrsbarOut_0_wordOffset1H,
  output [3:0] io_addrCrsbarOut_1_wordOffset1H,
  output [3:0] io_addrCrsbarOut_2_wordOffset1H,
  output [3:0] io_addrCrsbarOut_3_wordOffset1H,
  output [3:0] io_addrCrsbarOut_4_wordOffset1H,
  output [3:0] io_addrCrsbarOut_5_wordOffset1H,
  output [3:0] io_addrCrsbarOut_6_wordOffset1H,
  output [3:0] io_addrCrsbarOut_7_wordOffset1H,
  output       io_bankConflict
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  bankConflict_reg; // @[BankConflictArbiter.scala 103:33]
  reg  conflictReqIsW_reg; // @[BankConflictArbiter.scala 104:31]
  reg  perLaneConflictReq_reg_0_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_0_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_1_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_1_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_2_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_2_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_3_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_3_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_4_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_4_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_5_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_5_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_6_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_6_bankIdx; // @[BankConflictArbiter.scala 106:35]
  reg  perLaneConflictReq_reg_7_activeMask; // @[BankConflictArbiter.scala 106:35]
  reg [2:0] perLaneConflictReq_reg_7_bankIdx; // @[BankConflictArbiter.scala 106:35]
  wire  isWrite = bankConflict_reg ? conflictReqIsW_reg : io_coreReqArb_isWrite; // @[BankConflictArbiter.scala 121:26]
  wire [2:0] perLaneConflictReq_0_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_0_bankIdx :
    io_coreReqArb_perLaneAddr_0_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_0 = 8'h1 << perLaneConflictReq_0_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_0_activeMask = bankConflict_reg ? perLaneConflictReq_reg_0_activeMask :
    io_coreReqArb_perLaneAddr_0_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_0_T_1 = perLaneConflictReq_0_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_0 = bankIdx1H_0 & _bankIdxMasked_0_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_1_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_1_bankIdx :
    io_coreReqArb_perLaneAddr_1_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_1 = 8'h1 << perLaneConflictReq_1_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_1_activeMask = bankConflict_reg ? perLaneConflictReq_reg_1_activeMask :
    io_coreReqArb_perLaneAddr_1_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_1_T_1 = perLaneConflictReq_1_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_1 = bankIdx1H_1 & _bankIdxMasked_1_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_2_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_2_bankIdx :
    io_coreReqArb_perLaneAddr_2_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_2 = 8'h1 << perLaneConflictReq_2_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_2_activeMask = bankConflict_reg ? perLaneConflictReq_reg_2_activeMask :
    io_coreReqArb_perLaneAddr_2_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_2_T_1 = perLaneConflictReq_2_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_2 = bankIdx1H_2 & _bankIdxMasked_2_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_3_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_3_bankIdx :
    io_coreReqArb_perLaneAddr_3_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_3 = 8'h1 << perLaneConflictReq_3_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_3_activeMask = bankConflict_reg ? perLaneConflictReq_reg_3_activeMask :
    io_coreReqArb_perLaneAddr_3_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_3_T_1 = perLaneConflictReq_3_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_3 = bankIdx1H_3 & _bankIdxMasked_3_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_4_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_4_bankIdx :
    io_coreReqArb_perLaneAddr_4_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_4 = 8'h1 << perLaneConflictReq_4_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_4_activeMask = bankConflict_reg ? perLaneConflictReq_reg_4_activeMask :
    io_coreReqArb_perLaneAddr_4_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_4_T_1 = perLaneConflictReq_4_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_4 = bankIdx1H_4 & _bankIdxMasked_4_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_5_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_5_bankIdx :
    io_coreReqArb_perLaneAddr_5_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_5 = 8'h1 << perLaneConflictReq_5_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_5_activeMask = bankConflict_reg ? perLaneConflictReq_reg_5_activeMask :
    io_coreReqArb_perLaneAddr_5_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_5_T_1 = perLaneConflictReq_5_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_5 = bankIdx1H_5 & _bankIdxMasked_5_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_6_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_6_bankIdx :
    io_coreReqArb_perLaneAddr_6_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_6 = 8'h1 << perLaneConflictReq_6_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_6_activeMask = bankConflict_reg ? perLaneConflictReq_reg_6_activeMask :
    io_coreReqArb_perLaneAddr_6_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_6_T_1 = perLaneConflictReq_6_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_6 = bankIdx1H_6 & _bankIdxMasked_6_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [2:0] perLaneConflictReq_7_bankIdx = bankConflict_reg ? perLaneConflictReq_reg_7_bankIdx :
    io_coreReqArb_perLaneAddr_7_blockOffset; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] bankIdx1H_7 = 8'h1 << perLaneConflictReq_7_bankIdx; // @[OneHot.scala 57:35]
  wire  perLaneConflictReq_7_activeMask = bankConflict_reg ? perLaneConflictReq_reg_7_activeMask :
    io_coreReqArb_perLaneAddr_7_activeMask; // @[BankConflictArbiter.scala 157:28]
  wire [7:0] _bankIdxMasked_7_T_1 = perLaneConflictReq_7_activeMask ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] bankIdxMasked_7 = bankIdx1H_7 & _bankIdxMasked_7_T_1; // @[BankConflictArbiter.scala 129:38]
  wire [7:0] _perBankReq_Bin_0_T_8 = {bankIdxMasked_0[0],bankIdxMasked_1[0],bankIdxMasked_2[0],bankIdxMasked_3[0],
    bankIdxMasked_4[0],bankIdxMasked_5[0],bankIdxMasked_6[0],bankIdxMasked_7[0]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_17 = {{4'd0}, _perBankReq_Bin_0_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_12 = _GEN_17 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_14 = {_perBankReq_Bin_0_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_0_T_16 = _perBankReq_Bin_0_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_0_T_17 = _perBankReq_Bin_0_T_12 | _perBankReq_Bin_0_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_18 = {{2'd0}, _perBankReq_Bin_0_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_22 = _GEN_18 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_24 = {_perBankReq_Bin_0_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_0_T_26 = _perBankReq_Bin_0_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_0_T_27 = _perBankReq_Bin_0_T_22 | _perBankReq_Bin_0_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_19 = {{1'd0}, _perBankReq_Bin_0_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_32 = _GEN_19 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_0_T_34 = {_perBankReq_Bin_0_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_0_T_36 = _perBankReq_Bin_0_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_0 = _perBankReq_Bin_0_T_32 | _perBankReq_Bin_0_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_0_T_8 = perBankReq_Bin_0[0] + perBankReq_Bin_0[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_0_T_10 = perBankReq_Bin_0[2] + perBankReq_Bin_0[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_0_T_12 = _perBankReqCount_0_T_8 + _perBankReqCount_0_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_0_T_14 = perBankReq_Bin_0[4] + perBankReq_Bin_0[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_0_T_16 = perBankReq_Bin_0[6] + perBankReq_Bin_0[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_0_T_18 = _perBankReqCount_0_T_14 + _perBankReqCount_0_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_0_T_20 = _perBankReqCount_0_T_12 + _perBankReqCount_0_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_1_T_8 = {bankIdxMasked_0[1],bankIdxMasked_1[1],bankIdxMasked_2[1],bankIdxMasked_3[1],
    bankIdxMasked_4[1],bankIdxMasked_5[1],bankIdxMasked_6[1],bankIdxMasked_7[1]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_20 = {{4'd0}, _perBankReq_Bin_1_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_12 = _GEN_20 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_14 = {_perBankReq_Bin_1_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_1_T_16 = _perBankReq_Bin_1_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_1_T_17 = _perBankReq_Bin_1_T_12 | _perBankReq_Bin_1_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_21 = {{2'd0}, _perBankReq_Bin_1_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_22 = _GEN_21 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_24 = {_perBankReq_Bin_1_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_1_T_26 = _perBankReq_Bin_1_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_1_T_27 = _perBankReq_Bin_1_T_22 | _perBankReq_Bin_1_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_22 = {{1'd0}, _perBankReq_Bin_1_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_32 = _GEN_22 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_1_T_34 = {_perBankReq_Bin_1_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_1_T_36 = _perBankReq_Bin_1_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_1 = _perBankReq_Bin_1_T_32 | _perBankReq_Bin_1_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_1_T_8 = perBankReq_Bin_1[0] + perBankReq_Bin_1[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_1_T_10 = perBankReq_Bin_1[2] + perBankReq_Bin_1[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_1_T_12 = _perBankReqCount_1_T_8 + _perBankReqCount_1_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_1_T_14 = perBankReq_Bin_1[4] + perBankReq_Bin_1[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_1_T_16 = perBankReq_Bin_1[6] + perBankReq_Bin_1[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_1_T_18 = _perBankReqCount_1_T_14 + _perBankReqCount_1_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_1_T_20 = _perBankReqCount_1_T_12 + _perBankReqCount_1_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_2_T_8 = {bankIdxMasked_0[2],bankIdxMasked_1[2],bankIdxMasked_2[2],bankIdxMasked_3[2],
    bankIdxMasked_4[2],bankIdxMasked_5[2],bankIdxMasked_6[2],bankIdxMasked_7[2]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_23 = {{4'd0}, _perBankReq_Bin_2_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_12 = _GEN_23 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_14 = {_perBankReq_Bin_2_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_2_T_16 = _perBankReq_Bin_2_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_2_T_17 = _perBankReq_Bin_2_T_12 | _perBankReq_Bin_2_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_24 = {{2'd0}, _perBankReq_Bin_2_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_22 = _GEN_24 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_24 = {_perBankReq_Bin_2_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_2_T_26 = _perBankReq_Bin_2_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_2_T_27 = _perBankReq_Bin_2_T_22 | _perBankReq_Bin_2_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_25 = {{1'd0}, _perBankReq_Bin_2_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_32 = _GEN_25 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_2_T_34 = {_perBankReq_Bin_2_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_2_T_36 = _perBankReq_Bin_2_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_2 = _perBankReq_Bin_2_T_32 | _perBankReq_Bin_2_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_2_T_8 = perBankReq_Bin_2[0] + perBankReq_Bin_2[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_2_T_10 = perBankReq_Bin_2[2] + perBankReq_Bin_2[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_2_T_12 = _perBankReqCount_2_T_8 + _perBankReqCount_2_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_2_T_14 = perBankReq_Bin_2[4] + perBankReq_Bin_2[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_2_T_16 = perBankReq_Bin_2[6] + perBankReq_Bin_2[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_2_T_18 = _perBankReqCount_2_T_14 + _perBankReqCount_2_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_2_T_20 = _perBankReqCount_2_T_12 + _perBankReqCount_2_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_3_T_8 = {bankIdxMasked_0[3],bankIdxMasked_1[3],bankIdxMasked_2[3],bankIdxMasked_3[3],
    bankIdxMasked_4[3],bankIdxMasked_5[3],bankIdxMasked_6[3],bankIdxMasked_7[3]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_26 = {{4'd0}, _perBankReq_Bin_3_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_12 = _GEN_26 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_14 = {_perBankReq_Bin_3_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_3_T_16 = _perBankReq_Bin_3_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_3_T_17 = _perBankReq_Bin_3_T_12 | _perBankReq_Bin_3_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_27 = {{2'd0}, _perBankReq_Bin_3_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_22 = _GEN_27 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_24 = {_perBankReq_Bin_3_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_3_T_26 = _perBankReq_Bin_3_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_3_T_27 = _perBankReq_Bin_3_T_22 | _perBankReq_Bin_3_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_28 = {{1'd0}, _perBankReq_Bin_3_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_32 = _GEN_28 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_3_T_34 = {_perBankReq_Bin_3_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_3_T_36 = _perBankReq_Bin_3_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_3 = _perBankReq_Bin_3_T_32 | _perBankReq_Bin_3_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_3_T_8 = perBankReq_Bin_3[0] + perBankReq_Bin_3[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_3_T_10 = perBankReq_Bin_3[2] + perBankReq_Bin_3[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_3_T_12 = _perBankReqCount_3_T_8 + _perBankReqCount_3_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_3_T_14 = perBankReq_Bin_3[4] + perBankReq_Bin_3[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_3_T_16 = perBankReq_Bin_3[6] + perBankReq_Bin_3[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_3_T_18 = _perBankReqCount_3_T_14 + _perBankReqCount_3_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_3_T_20 = _perBankReqCount_3_T_12 + _perBankReqCount_3_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_4_T_8 = {bankIdxMasked_0[4],bankIdxMasked_1[4],bankIdxMasked_2[4],bankIdxMasked_3[4],
    bankIdxMasked_4[4],bankIdxMasked_5[4],bankIdxMasked_6[4],bankIdxMasked_7[4]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_29 = {{4'd0}, _perBankReq_Bin_4_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_12 = _GEN_29 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_14 = {_perBankReq_Bin_4_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_4_T_16 = _perBankReq_Bin_4_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_4_T_17 = _perBankReq_Bin_4_T_12 | _perBankReq_Bin_4_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_30 = {{2'd0}, _perBankReq_Bin_4_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_22 = _GEN_30 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_24 = {_perBankReq_Bin_4_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_4_T_26 = _perBankReq_Bin_4_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_4_T_27 = _perBankReq_Bin_4_T_22 | _perBankReq_Bin_4_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_31 = {{1'd0}, _perBankReq_Bin_4_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_32 = _GEN_31 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_4_T_34 = {_perBankReq_Bin_4_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_4_T_36 = _perBankReq_Bin_4_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_4 = _perBankReq_Bin_4_T_32 | _perBankReq_Bin_4_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_4_T_8 = perBankReq_Bin_4[0] + perBankReq_Bin_4[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_4_T_10 = perBankReq_Bin_4[2] + perBankReq_Bin_4[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_4_T_12 = _perBankReqCount_4_T_8 + _perBankReqCount_4_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_4_T_14 = perBankReq_Bin_4[4] + perBankReq_Bin_4[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_4_T_16 = perBankReq_Bin_4[6] + perBankReq_Bin_4[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_4_T_18 = _perBankReqCount_4_T_14 + _perBankReqCount_4_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_4_T_20 = _perBankReqCount_4_T_12 + _perBankReqCount_4_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_5_T_8 = {bankIdxMasked_0[5],bankIdxMasked_1[5],bankIdxMasked_2[5],bankIdxMasked_3[5],
    bankIdxMasked_4[5],bankIdxMasked_5[5],bankIdxMasked_6[5],bankIdxMasked_7[5]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_32 = {{4'd0}, _perBankReq_Bin_5_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_12 = _GEN_32 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_14 = {_perBankReq_Bin_5_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_5_T_16 = _perBankReq_Bin_5_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_5_T_17 = _perBankReq_Bin_5_T_12 | _perBankReq_Bin_5_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_33 = {{2'd0}, _perBankReq_Bin_5_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_22 = _GEN_33 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_24 = {_perBankReq_Bin_5_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_5_T_26 = _perBankReq_Bin_5_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_5_T_27 = _perBankReq_Bin_5_T_22 | _perBankReq_Bin_5_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_34 = {{1'd0}, _perBankReq_Bin_5_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_32 = _GEN_34 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_5_T_34 = {_perBankReq_Bin_5_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_5_T_36 = _perBankReq_Bin_5_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_5 = _perBankReq_Bin_5_T_32 | _perBankReq_Bin_5_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_5_T_8 = perBankReq_Bin_5[0] + perBankReq_Bin_5[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_5_T_10 = perBankReq_Bin_5[2] + perBankReq_Bin_5[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_5_T_12 = _perBankReqCount_5_T_8 + _perBankReqCount_5_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_5_T_14 = perBankReq_Bin_5[4] + perBankReq_Bin_5[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_5_T_16 = perBankReq_Bin_5[6] + perBankReq_Bin_5[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_5_T_18 = _perBankReqCount_5_T_14 + _perBankReqCount_5_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_5_T_20 = _perBankReqCount_5_T_12 + _perBankReqCount_5_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_6_T_8 = {bankIdxMasked_0[6],bankIdxMasked_1[6],bankIdxMasked_2[6],bankIdxMasked_3[6],
    bankIdxMasked_4[6],bankIdxMasked_5[6],bankIdxMasked_6[6],bankIdxMasked_7[6]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_35 = {{4'd0}, _perBankReq_Bin_6_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_12 = _GEN_35 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_14 = {_perBankReq_Bin_6_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_6_T_16 = _perBankReq_Bin_6_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_6_T_17 = _perBankReq_Bin_6_T_12 | _perBankReq_Bin_6_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_36 = {{2'd0}, _perBankReq_Bin_6_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_22 = _GEN_36 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_24 = {_perBankReq_Bin_6_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_6_T_26 = _perBankReq_Bin_6_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_6_T_27 = _perBankReq_Bin_6_T_22 | _perBankReq_Bin_6_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_37 = {{1'd0}, _perBankReq_Bin_6_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_32 = _GEN_37 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_6_T_34 = {_perBankReq_Bin_6_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_6_T_36 = _perBankReq_Bin_6_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_6 = _perBankReq_Bin_6_T_32 | _perBankReq_Bin_6_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_6_T_8 = perBankReq_Bin_6[0] + perBankReq_Bin_6[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_6_T_10 = perBankReq_Bin_6[2] + perBankReq_Bin_6[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_6_T_12 = _perBankReqCount_6_T_8 + _perBankReqCount_6_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_6_T_14 = perBankReq_Bin_6[4] + perBankReq_Bin_6[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_6_T_16 = perBankReq_Bin_6[6] + perBankReq_Bin_6[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_6_T_18 = _perBankReqCount_6_T_14 + _perBankReqCount_6_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_6_T_20 = _perBankReqCount_6_T_12 + _perBankReqCount_6_T_18; // @[Bitwise.scala 48:55]
  wire [7:0] _perBankReq_Bin_7_T_8 = {bankIdxMasked_0[7],bankIdxMasked_1[7],bankIdxMasked_2[7],bankIdxMasked_3[7],
    bankIdxMasked_4[7],bankIdxMasked_5[7],bankIdxMasked_6[7],bankIdxMasked_7[7]}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_38 = {{4'd0}, _perBankReq_Bin_7_T_8[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_12 = _GEN_38 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_14 = {_perBankReq_Bin_7_T_8[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_7_T_16 = _perBankReq_Bin_7_T_14 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_7_T_17 = _perBankReq_Bin_7_T_12 | _perBankReq_Bin_7_T_16; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_39 = {{2'd0}, _perBankReq_Bin_7_T_17[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_22 = _GEN_39 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_24 = {_perBankReq_Bin_7_T_17[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_7_T_26 = _perBankReq_Bin_7_T_24 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _perBankReq_Bin_7_T_27 = _perBankReq_Bin_7_T_22 | _perBankReq_Bin_7_T_26; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_40 = {{1'd0}, _perBankReq_Bin_7_T_27[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_32 = _GEN_40 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _perBankReq_Bin_7_T_34 = {_perBankReq_Bin_7_T_27[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _perBankReq_Bin_7_T_36 = _perBankReq_Bin_7_T_34 & 8'haa; // @[Bitwise.scala 105:80]
  wire [7:0] perBankReq_Bin_7 = _perBankReq_Bin_7_T_32 | _perBankReq_Bin_7_T_36; // @[Bitwise.scala 105:39]
  wire [1:0] _perBankReqCount_7_T_8 = perBankReq_Bin_7[0] + perBankReq_Bin_7[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_7_T_10 = perBankReq_Bin_7[2] + perBankReq_Bin_7[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_7_T_12 = _perBankReqCount_7_T_8 + _perBankReqCount_7_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_7_T_14 = perBankReq_Bin_7[4] + perBankReq_Bin_7[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _perBankReqCount_7_T_16 = perBankReq_Bin_7[6] + perBankReq_Bin_7[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _perBankReqCount_7_T_18 = _perBankReqCount_7_T_14 + _perBankReqCount_7_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _perBankReqCount_7_T_20 = _perBankReqCount_7_T_12 + _perBankReqCount_7_T_18; // @[Bitwise.scala 48:55]
  wire [2:0] perBankReqCount_0 = _perBankReqCount_0_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_0 = perBankReqCount_0 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_1 = _perBankReqCount_1_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_1 = perBankReqCount_1 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_2 = _perBankReqCount_2_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_2 = perBankReqCount_2 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_3 = _perBankReqCount_3_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_3 = perBankReqCount_3 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_4 = _perBankReqCount_4_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_4 = perBankReqCount_4 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_5 = _perBankReqCount_5_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_5 = perBankReqCount_5 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_6 = _perBankReqCount_6_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_6 = perBankReqCount_6 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [2:0] perBankReqCount_7 = _perBankReqCount_7_T_20[2:0]; // @[BankConflictArbiter.scala 131:29 134:24]
  wire  perBankReqConflict_7 = perBankReqCount_7 > 3'h1; // @[BankConflictArbiter.scala 145:46]
  wire [7:0] _bankConflict_T = {perBankReqConflict_0,perBankReqConflict_1,perBankReqConflict_2,perBankReqConflict_3,
    perBankReqConflict_4,perBankReqConflict_5,perBankReqConflict_6,perBankReqConflict_7}; // @[Cat.scala 31:58]
  wire  bankConflict = |_bankConflict_T; // @[BankConflictArbiter.scala 146:43]
  wire [7:0] _T_16 = perBankReq_Bin_0[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_17 = perBankReq_Bin_0[6] ? 8'h40 : _T_16; // @[Mux.scala 47:70]
  wire [7:0] _T_18 = perBankReq_Bin_0[5] ? 8'h20 : _T_17; // @[Mux.scala 47:70]
  wire [7:0] _T_19 = perBankReq_Bin_0[4] ? 8'h10 : _T_18; // @[Mux.scala 47:70]
  wire [7:0] _T_20 = perBankReq_Bin_0[3] ? 8'h8 : _T_19; // @[Mux.scala 47:70]
  wire [7:0] _T_21 = perBankReq_Bin_0[2] ? 8'h4 : _T_20; // @[Mux.scala 47:70]
  wire [7:0] _T_22 = perBankReq_Bin_0[1] ? 8'h2 : _T_21; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_0 = perBankReq_Bin_0[0] ? 8'h1 : _T_22; // @[Mux.scala 47:70]
  wire [7:0] _T_32 = perBankReq_Bin_1[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_33 = perBankReq_Bin_1[6] ? 8'h40 : _T_32; // @[Mux.scala 47:70]
  wire [7:0] _T_34 = perBankReq_Bin_1[5] ? 8'h20 : _T_33; // @[Mux.scala 47:70]
  wire [7:0] _T_35 = perBankReq_Bin_1[4] ? 8'h10 : _T_34; // @[Mux.scala 47:70]
  wire [7:0] _T_36 = perBankReq_Bin_1[3] ? 8'h8 : _T_35; // @[Mux.scala 47:70]
  wire [7:0] _T_37 = perBankReq_Bin_1[2] ? 8'h4 : _T_36; // @[Mux.scala 47:70]
  wire [7:0] _T_38 = perBankReq_Bin_1[1] ? 8'h2 : _T_37; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_1 = perBankReq_Bin_1[0] ? 8'h1 : _T_38; // @[Mux.scala 47:70]
  wire [7:0] _T_48 = perBankReq_Bin_2[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_49 = perBankReq_Bin_2[6] ? 8'h40 : _T_48; // @[Mux.scala 47:70]
  wire [7:0] _T_50 = perBankReq_Bin_2[5] ? 8'h20 : _T_49; // @[Mux.scala 47:70]
  wire [7:0] _T_51 = perBankReq_Bin_2[4] ? 8'h10 : _T_50; // @[Mux.scala 47:70]
  wire [7:0] _T_52 = perBankReq_Bin_2[3] ? 8'h8 : _T_51; // @[Mux.scala 47:70]
  wire [7:0] _T_53 = perBankReq_Bin_2[2] ? 8'h4 : _T_52; // @[Mux.scala 47:70]
  wire [7:0] _T_54 = perBankReq_Bin_2[1] ? 8'h2 : _T_53; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_2 = perBankReq_Bin_2[0] ? 8'h1 : _T_54; // @[Mux.scala 47:70]
  wire [7:0] _T_64 = perBankReq_Bin_3[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_65 = perBankReq_Bin_3[6] ? 8'h40 : _T_64; // @[Mux.scala 47:70]
  wire [7:0] _T_66 = perBankReq_Bin_3[5] ? 8'h20 : _T_65; // @[Mux.scala 47:70]
  wire [7:0] _T_67 = perBankReq_Bin_3[4] ? 8'h10 : _T_66; // @[Mux.scala 47:70]
  wire [7:0] _T_68 = perBankReq_Bin_3[3] ? 8'h8 : _T_67; // @[Mux.scala 47:70]
  wire [7:0] _T_69 = perBankReq_Bin_3[2] ? 8'h4 : _T_68; // @[Mux.scala 47:70]
  wire [7:0] _T_70 = perBankReq_Bin_3[1] ? 8'h2 : _T_69; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_3 = perBankReq_Bin_3[0] ? 8'h1 : _T_70; // @[Mux.scala 47:70]
  wire [7:0] _T_80 = perBankReq_Bin_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_81 = perBankReq_Bin_4[6] ? 8'h40 : _T_80; // @[Mux.scala 47:70]
  wire [7:0] _T_82 = perBankReq_Bin_4[5] ? 8'h20 : _T_81; // @[Mux.scala 47:70]
  wire [7:0] _T_83 = perBankReq_Bin_4[4] ? 8'h10 : _T_82; // @[Mux.scala 47:70]
  wire [7:0] _T_84 = perBankReq_Bin_4[3] ? 8'h8 : _T_83; // @[Mux.scala 47:70]
  wire [7:0] _T_85 = perBankReq_Bin_4[2] ? 8'h4 : _T_84; // @[Mux.scala 47:70]
  wire [7:0] _T_86 = perBankReq_Bin_4[1] ? 8'h2 : _T_85; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_4 = perBankReq_Bin_4[0] ? 8'h1 : _T_86; // @[Mux.scala 47:70]
  wire [7:0] _T_96 = perBankReq_Bin_5[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_97 = perBankReq_Bin_5[6] ? 8'h40 : _T_96; // @[Mux.scala 47:70]
  wire [7:0] _T_98 = perBankReq_Bin_5[5] ? 8'h20 : _T_97; // @[Mux.scala 47:70]
  wire [7:0] _T_99 = perBankReq_Bin_5[4] ? 8'h10 : _T_98; // @[Mux.scala 47:70]
  wire [7:0] _T_100 = perBankReq_Bin_5[3] ? 8'h8 : _T_99; // @[Mux.scala 47:70]
  wire [7:0] _T_101 = perBankReq_Bin_5[2] ? 8'h4 : _T_100; // @[Mux.scala 47:70]
  wire [7:0] _T_102 = perBankReq_Bin_5[1] ? 8'h2 : _T_101; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_5 = perBankReq_Bin_5[0] ? 8'h1 : _T_102; // @[Mux.scala 47:70]
  wire [7:0] _T_112 = perBankReq_Bin_6[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_113 = perBankReq_Bin_6[6] ? 8'h40 : _T_112; // @[Mux.scala 47:70]
  wire [7:0] _T_114 = perBankReq_Bin_6[5] ? 8'h20 : _T_113; // @[Mux.scala 47:70]
  wire [7:0] _T_115 = perBankReq_Bin_6[4] ? 8'h10 : _T_114; // @[Mux.scala 47:70]
  wire [7:0] _T_116 = perBankReq_Bin_6[3] ? 8'h8 : _T_115; // @[Mux.scala 47:70]
  wire [7:0] _T_117 = perBankReq_Bin_6[2] ? 8'h4 : _T_116; // @[Mux.scala 47:70]
  wire [7:0] _T_118 = perBankReq_Bin_6[1] ? 8'h2 : _T_117; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_6 = perBankReq_Bin_6[0] ? 8'h1 : _T_118; // @[Mux.scala 47:70]
  wire [7:0] _T_128 = perBankReq_Bin_7[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _T_129 = perBankReq_Bin_7[6] ? 8'h40 : _T_128; // @[Mux.scala 47:70]
  wire [7:0] _T_130 = perBankReq_Bin_7[5] ? 8'h20 : _T_129; // @[Mux.scala 47:70]
  wire [7:0] _T_131 = perBankReq_Bin_7[4] ? 8'h10 : _T_130; // @[Mux.scala 47:70]
  wire [7:0] _T_132 = perBankReq_Bin_7[3] ? 8'h8 : _T_131; // @[Mux.scala 47:70]
  wire [7:0] _T_133 = perBankReq_Bin_7[2] ? 8'h4 : _T_132; // @[Mux.scala 47:70]
  wire [7:0] _T_134 = perBankReq_Bin_7[1] ? 8'h2 : _T_133; // @[Mux.scala 47:70]
  wire [7:0] perBankActiveLaneWhenConflict1H_7 = perBankReq_Bin_7[0] ? 8'h1 : _T_134; // @[Mux.scala 47:70]
  wire [7:0] _ActiveLaneWhenConflict1H_0_T_8 = {perBankActiveLaneWhenConflict1H_0[0],perBankActiveLaneWhenConflict1H_1[0
    ],perBankActiveLaneWhenConflict1H_2[0],perBankActiveLaneWhenConflict1H_3[0],perBankActiveLaneWhenConflict1H_4[0],
    perBankActiveLaneWhenConflict1H_5[0],perBankActiveLaneWhenConflict1H_6[0],perBankActiveLaneWhenConflict1H_7[0]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_0 = |_ActiveLaneWhenConflict1H_0_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_1_T_8 = {perBankActiveLaneWhenConflict1H_0[1],perBankActiveLaneWhenConflict1H_1[1
    ],perBankActiveLaneWhenConflict1H_2[1],perBankActiveLaneWhenConflict1H_3[1],perBankActiveLaneWhenConflict1H_4[1],
    perBankActiveLaneWhenConflict1H_5[1],perBankActiveLaneWhenConflict1H_6[1],perBankActiveLaneWhenConflict1H_7[1]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_1 = |_ActiveLaneWhenConflict1H_1_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_2_T_8 = {perBankActiveLaneWhenConflict1H_0[2],perBankActiveLaneWhenConflict1H_1[2
    ],perBankActiveLaneWhenConflict1H_2[2],perBankActiveLaneWhenConflict1H_3[2],perBankActiveLaneWhenConflict1H_4[2],
    perBankActiveLaneWhenConflict1H_5[2],perBankActiveLaneWhenConflict1H_6[2],perBankActiveLaneWhenConflict1H_7[2]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_2 = |_ActiveLaneWhenConflict1H_2_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_3_T_8 = {perBankActiveLaneWhenConflict1H_0[3],perBankActiveLaneWhenConflict1H_1[3
    ],perBankActiveLaneWhenConflict1H_2[3],perBankActiveLaneWhenConflict1H_3[3],perBankActiveLaneWhenConflict1H_4[3],
    perBankActiveLaneWhenConflict1H_5[3],perBankActiveLaneWhenConflict1H_6[3],perBankActiveLaneWhenConflict1H_7[3]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_3 = |_ActiveLaneWhenConflict1H_3_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_4_T_8 = {perBankActiveLaneWhenConflict1H_0[4],perBankActiveLaneWhenConflict1H_1[4
    ],perBankActiveLaneWhenConflict1H_2[4],perBankActiveLaneWhenConflict1H_3[4],perBankActiveLaneWhenConflict1H_4[4],
    perBankActiveLaneWhenConflict1H_5[4],perBankActiveLaneWhenConflict1H_6[4],perBankActiveLaneWhenConflict1H_7[4]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_4 = |_ActiveLaneWhenConflict1H_4_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_5_T_8 = {perBankActiveLaneWhenConflict1H_0[5],perBankActiveLaneWhenConflict1H_1[5
    ],perBankActiveLaneWhenConflict1H_2[5],perBankActiveLaneWhenConflict1H_3[5],perBankActiveLaneWhenConflict1H_4[5],
    perBankActiveLaneWhenConflict1H_5[5],perBankActiveLaneWhenConflict1H_6[5],perBankActiveLaneWhenConflict1H_7[5]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_5 = |_ActiveLaneWhenConflict1H_5_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_6_T_8 = {perBankActiveLaneWhenConflict1H_0[6],perBankActiveLaneWhenConflict1H_1[6
    ],perBankActiveLaneWhenConflict1H_2[6],perBankActiveLaneWhenConflict1H_3[6],perBankActiveLaneWhenConflict1H_4[6],
    perBankActiveLaneWhenConflict1H_5[6],perBankActiveLaneWhenConflict1H_6[6],perBankActiveLaneWhenConflict1H_7[6]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_6 = |_ActiveLaneWhenConflict1H_6_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ActiveLaneWhenConflict1H_7_T_8 = {perBankActiveLaneWhenConflict1H_0[7],perBankActiveLaneWhenConflict1H_1[7
    ],perBankActiveLaneWhenConflict1H_2[7],perBankActiveLaneWhenConflict1H_3[7],perBankActiveLaneWhenConflict1H_4[7],
    perBankActiveLaneWhenConflict1H_5[7],perBankActiveLaneWhenConflict1H_6[7],perBankActiveLaneWhenConflict1H_7[7]}; // @[Cat.scala 31:58]
  wire  ActiveLaneWhenConflict1H_7 = |_ActiveLaneWhenConflict1H_7_T_8; // @[BankConflictArbiter.scala 154:83]
  wire [7:0] _ReserveLaneWhenConflict1H_T = {ActiveLaneWhenConflict1H_0,ActiveLaneWhenConflict1H_1,
    ActiveLaneWhenConflict1H_2,ActiveLaneWhenConflict1H_3,ActiveLaneWhenConflict1H_4,ActiveLaneWhenConflict1H_5,
    ActiveLaneWhenConflict1H_6,ActiveLaneWhenConflict1H_7}; // @[Cat.scala 31:58]
  wire [7:0] _ReserveLaneWhenConflict1H_T_1 = {perLaneConflictReq_0_activeMask,perLaneConflictReq_1_activeMask,
    perLaneConflictReq_2_activeMask,perLaneConflictReq_3_activeMask,perLaneConflictReq_4_activeMask,
    perLaneConflictReq_5_activeMask,perLaneConflictReq_6_activeMask,perLaneConflictReq_7_activeMask}; // @[Cat.scala 31:58]
  wire [7:0] _ReserveLaneWhenConflict1H_T_2 = _ReserveLaneWhenConflict1H_T & _ReserveLaneWhenConflict1H_T_1; // @[BankConflictArbiter.scala 155:74]
  wire  ReserveLaneWhenConflict1H_0 = _ReserveLaneWhenConflict1H_T_2[0]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_1 = _ReserveLaneWhenConflict1H_T_2[1]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_2 = _ReserveLaneWhenConflict1H_T_2[2]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_3 = _ReserveLaneWhenConflict1H_T_2[3]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_4 = _ReserveLaneWhenConflict1H_T_2[4]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_5 = _ReserveLaneWhenConflict1H_T_2[5]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_6 = _ReserveLaneWhenConflict1H_T_2[6]; // @[BankConflictArbiter.scala 155:97]
  wire  ReserveLaneWhenConflict1H_7 = _ReserveLaneWhenConflict1H_T_2[7]; // @[BankConflictArbiter.scala 155:97]
  wire [3:0] _T_145 = perBankActiveLaneWhenConflict1H_0[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_146 = perBankActiveLaneWhenConflict1H_0[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_147 = perBankActiveLaneWhenConflict1H_0[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_148 = perBankActiveLaneWhenConflict1H_0[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_149 = perBankActiveLaneWhenConflict1H_0[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_150 = perBankActiveLaneWhenConflict1H_0[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_151 = perBankActiveLaneWhenConflict1H_0[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_152 = perBankActiveLaneWhenConflict1H_0[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_153 = _T_145 | _T_146; // @[Mux.scala 27:73]
  wire [3:0] _T_154 = _T_153 | _T_147; // @[Mux.scala 27:73]
  wire [3:0] _T_155 = _T_154 | _T_148; // @[Mux.scala 27:73]
  wire [3:0] _T_156 = _T_155 | _T_149; // @[Mux.scala 27:73]
  wire [3:0] _T_157 = _T_156 | _T_150; // @[Mux.scala 27:73]
  wire [3:0] _T_158 = _T_157 | _T_151; // @[Mux.scala 27:73]
  wire [3:0] _T_168 = perBankActiveLaneWhenConflict1H_1[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_169 = perBankActiveLaneWhenConflict1H_1[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_170 = perBankActiveLaneWhenConflict1H_1[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_171 = perBankActiveLaneWhenConflict1H_1[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_172 = perBankActiveLaneWhenConflict1H_1[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_173 = perBankActiveLaneWhenConflict1H_1[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_174 = perBankActiveLaneWhenConflict1H_1[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_175 = perBankActiveLaneWhenConflict1H_1[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_176 = _T_168 | _T_169; // @[Mux.scala 27:73]
  wire [3:0] _T_177 = _T_176 | _T_170; // @[Mux.scala 27:73]
  wire [3:0] _T_178 = _T_177 | _T_171; // @[Mux.scala 27:73]
  wire [3:0] _T_179 = _T_178 | _T_172; // @[Mux.scala 27:73]
  wire [3:0] _T_180 = _T_179 | _T_173; // @[Mux.scala 27:73]
  wire [3:0] _T_181 = _T_180 | _T_174; // @[Mux.scala 27:73]
  wire [3:0] _T_191 = perBankActiveLaneWhenConflict1H_2[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_192 = perBankActiveLaneWhenConflict1H_2[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_193 = perBankActiveLaneWhenConflict1H_2[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_194 = perBankActiveLaneWhenConflict1H_2[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_195 = perBankActiveLaneWhenConflict1H_2[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_196 = perBankActiveLaneWhenConflict1H_2[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_197 = perBankActiveLaneWhenConflict1H_2[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_198 = perBankActiveLaneWhenConflict1H_2[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_199 = _T_191 | _T_192; // @[Mux.scala 27:73]
  wire [3:0] _T_200 = _T_199 | _T_193; // @[Mux.scala 27:73]
  wire [3:0] _T_201 = _T_200 | _T_194; // @[Mux.scala 27:73]
  wire [3:0] _T_202 = _T_201 | _T_195; // @[Mux.scala 27:73]
  wire [3:0] _T_203 = _T_202 | _T_196; // @[Mux.scala 27:73]
  wire [3:0] _T_204 = _T_203 | _T_197; // @[Mux.scala 27:73]
  wire [3:0] _T_214 = perBankActiveLaneWhenConflict1H_3[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_215 = perBankActiveLaneWhenConflict1H_3[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_216 = perBankActiveLaneWhenConflict1H_3[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_217 = perBankActiveLaneWhenConflict1H_3[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_218 = perBankActiveLaneWhenConflict1H_3[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_219 = perBankActiveLaneWhenConflict1H_3[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_220 = perBankActiveLaneWhenConflict1H_3[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_221 = perBankActiveLaneWhenConflict1H_3[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_222 = _T_214 | _T_215; // @[Mux.scala 27:73]
  wire [3:0] _T_223 = _T_222 | _T_216; // @[Mux.scala 27:73]
  wire [3:0] _T_224 = _T_223 | _T_217; // @[Mux.scala 27:73]
  wire [3:0] _T_225 = _T_224 | _T_218; // @[Mux.scala 27:73]
  wire [3:0] _T_226 = _T_225 | _T_219; // @[Mux.scala 27:73]
  wire [3:0] _T_227 = _T_226 | _T_220; // @[Mux.scala 27:73]
  wire [3:0] _T_237 = perBankActiveLaneWhenConflict1H_4[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_238 = perBankActiveLaneWhenConflict1H_4[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_239 = perBankActiveLaneWhenConflict1H_4[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_240 = perBankActiveLaneWhenConflict1H_4[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_241 = perBankActiveLaneWhenConflict1H_4[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_242 = perBankActiveLaneWhenConflict1H_4[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_243 = perBankActiveLaneWhenConflict1H_4[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_244 = perBankActiveLaneWhenConflict1H_4[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_245 = _T_237 | _T_238; // @[Mux.scala 27:73]
  wire [3:0] _T_246 = _T_245 | _T_239; // @[Mux.scala 27:73]
  wire [3:0] _T_247 = _T_246 | _T_240; // @[Mux.scala 27:73]
  wire [3:0] _T_248 = _T_247 | _T_241; // @[Mux.scala 27:73]
  wire [3:0] _T_249 = _T_248 | _T_242; // @[Mux.scala 27:73]
  wire [3:0] _T_250 = _T_249 | _T_243; // @[Mux.scala 27:73]
  wire [3:0] _T_260 = perBankActiveLaneWhenConflict1H_5[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_261 = perBankActiveLaneWhenConflict1H_5[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_262 = perBankActiveLaneWhenConflict1H_5[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_263 = perBankActiveLaneWhenConflict1H_5[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_264 = perBankActiveLaneWhenConflict1H_5[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_265 = perBankActiveLaneWhenConflict1H_5[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_266 = perBankActiveLaneWhenConflict1H_5[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_267 = perBankActiveLaneWhenConflict1H_5[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_268 = _T_260 | _T_261; // @[Mux.scala 27:73]
  wire [3:0] _T_269 = _T_268 | _T_262; // @[Mux.scala 27:73]
  wire [3:0] _T_270 = _T_269 | _T_263; // @[Mux.scala 27:73]
  wire [3:0] _T_271 = _T_270 | _T_264; // @[Mux.scala 27:73]
  wire [3:0] _T_272 = _T_271 | _T_265; // @[Mux.scala 27:73]
  wire [3:0] _T_273 = _T_272 | _T_266; // @[Mux.scala 27:73]
  wire [3:0] _T_283 = perBankActiveLaneWhenConflict1H_6[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_284 = perBankActiveLaneWhenConflict1H_6[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_285 = perBankActiveLaneWhenConflict1H_6[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_286 = perBankActiveLaneWhenConflict1H_6[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_287 = perBankActiveLaneWhenConflict1H_6[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_288 = perBankActiveLaneWhenConflict1H_6[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_289 = perBankActiveLaneWhenConflict1H_6[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_290 = perBankActiveLaneWhenConflict1H_6[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_291 = _T_283 | _T_284; // @[Mux.scala 27:73]
  wire [3:0] _T_292 = _T_291 | _T_285; // @[Mux.scala 27:73]
  wire [3:0] _T_293 = _T_292 | _T_286; // @[Mux.scala 27:73]
  wire [3:0] _T_294 = _T_293 | _T_287; // @[Mux.scala 27:73]
  wire [3:0] _T_295 = _T_294 | _T_288; // @[Mux.scala 27:73]
  wire [3:0] _T_296 = _T_295 | _T_289; // @[Mux.scala 27:73]
  wire [3:0] _T_306 = perBankActiveLaneWhenConflict1H_7[0] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_307 = perBankActiveLaneWhenConflict1H_7[1] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_308 = perBankActiveLaneWhenConflict1H_7[2] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_309 = perBankActiveLaneWhenConflict1H_7[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_310 = perBankActiveLaneWhenConflict1H_7[4] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_311 = perBankActiveLaneWhenConflict1H_7[5] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_312 = perBankActiveLaneWhenConflict1H_7[6] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_313 = perBankActiveLaneWhenConflict1H_7[7] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_314 = _T_306 | _T_307; // @[Mux.scala 27:73]
  wire [3:0] _T_315 = _T_314 | _T_308; // @[Mux.scala 27:73]
  wire [3:0] _T_316 = _T_315 | _T_309; // @[Mux.scala 27:73]
  wire [3:0] _T_317 = _T_316 | _T_310; // @[Mux.scala 27:73]
  wire [3:0] _T_318 = _T_317 | _T_311; // @[Mux.scala 27:73]
  wire [3:0] _T_319 = _T_318 | _T_312; // @[Mux.scala 27:73]
  assign io_dataCrsbarSel1H_0 = isWrite ? perBankActiveLaneWhenConflict1H_0 : bankIdxMasked_0; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_1 = isWrite ? perBankActiveLaneWhenConflict1H_1 : bankIdxMasked_1; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_2 = isWrite ? perBankActiveLaneWhenConflict1H_2 : bankIdxMasked_2; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_3 = isWrite ? perBankActiveLaneWhenConflict1H_3 : bankIdxMasked_3; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_4 = isWrite ? perBankActiveLaneWhenConflict1H_4 : bankIdxMasked_4; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_5 = isWrite ? perBankActiveLaneWhenConflict1H_5 : bankIdxMasked_5; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_6 = isWrite ? perBankActiveLaneWhenConflict1H_6 : bankIdxMasked_6; // @[BankConflictArbiter.scala 172:28]
  assign io_dataCrsbarSel1H_7 = isWrite ? perBankActiveLaneWhenConflict1H_7 : bankIdxMasked_7; // @[BankConflictArbiter.scala 172:28]
  assign io_addrCrsbarOut_0_wordOffset1H = _T_158 | _T_152; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_1_wordOffset1H = _T_181 | _T_175; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_2_wordOffset1H = _T_204 | _T_198; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_3_wordOffset1H = _T_227 | _T_221; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_4_wordOffset1H = _T_250 | _T_244; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_5_wordOffset1H = _T_273 | _T_267; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_6_wordOffset1H = _T_296 | _T_290; // @[Mux.scala 27:73]
  assign io_addrCrsbarOut_7_wordOffset1H = _T_319 | _T_313; // @[Mux.scala 27:73]
  assign io_bankConflict = |_bankConflict_T; // @[BankConflictArbiter.scala 146:43]
  always @(posedge clock) begin
    if (reset) begin // @[BankConflictArbiter.scala 103:33]
      bankConflict_reg <= 1'h0; // @[BankConflictArbiter.scala 103:33]
    end else begin
      bankConflict_reg <= bankConflict; // @[BankConflictArbiter.scala 103:33]
    end
    if (bankConflict) begin // @[BankConflictArbiter.scala 165:21]
      conflictReqIsW_reg <= io_coreReqArb_isWrite; // @[BankConflictArbiter.scala 165:41]
    end
    perLaneConflictReq_reg_0_activeMask <= _ReserveLaneWhenConflict1H_T_2[0]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_0) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_0_bankIdx <= io_coreReqArb_perLaneAddr_0_blockOffset;
      end
    end
    perLaneConflictReq_reg_1_activeMask <= _ReserveLaneWhenConflict1H_T_2[1]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_1) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_1_bankIdx <= io_coreReqArb_perLaneAddr_1_blockOffset;
      end
    end
    perLaneConflictReq_reg_2_activeMask <= _ReserveLaneWhenConflict1H_T_2[2]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_2) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_2_bankIdx <= io_coreReqArb_perLaneAddr_2_blockOffset;
      end
    end
    perLaneConflictReq_reg_3_activeMask <= _ReserveLaneWhenConflict1H_T_2[3]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_3) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_3_bankIdx <= io_coreReqArb_perLaneAddr_3_blockOffset;
      end
    end
    perLaneConflictReq_reg_4_activeMask <= _ReserveLaneWhenConflict1H_T_2[4]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_4) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_4_bankIdx <= io_coreReqArb_perLaneAddr_4_blockOffset;
      end
    end
    perLaneConflictReq_reg_5_activeMask <= _ReserveLaneWhenConflict1H_T_2[5]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_5) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_5_bankIdx <= io_coreReqArb_perLaneAddr_5_blockOffset;
      end
    end
    perLaneConflictReq_reg_6_activeMask <= _ReserveLaneWhenConflict1H_T_2[6]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_6) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_6_bankIdx <= io_coreReqArb_perLaneAddr_6_blockOffset;
      end
    end
    perLaneConflictReq_reg_7_activeMask <= _ReserveLaneWhenConflict1H_T_2[7]; // @[BankConflictArbiter.scala 155:97]
    if (ReserveLaneWhenConflict1H_7) begin // @[BankConflictArbiter.scala 160:39]
      if (!(bankConflict_reg)) begin // @[BankConflictArbiter.scala 157:28]
        perLaneConflictReq_reg_7_bankIdx <= io_coreReqArb_perLaneAddr_7_blockOffset;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bankConflict_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  conflictReqIsW_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  perLaneConflictReq_reg_0_activeMask = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  perLaneConflictReq_reg_0_bankIdx = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  perLaneConflictReq_reg_1_activeMask = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  perLaneConflictReq_reg_1_bankIdx = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  perLaneConflictReq_reg_2_activeMask = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  perLaneConflictReq_reg_2_bankIdx = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  perLaneConflictReq_reg_3_activeMask = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  perLaneConflictReq_reg_3_bankIdx = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  perLaneConflictReq_reg_4_activeMask = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  perLaneConflictReq_reg_4_bankIdx = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  perLaneConflictReq_reg_5_activeMask = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  perLaneConflictReq_reg_5_bankIdx = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  perLaneConflictReq_reg_6_activeMask = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  perLaneConflictReq_reg_6_bankIdx = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  perLaneConflictReq_reg_7_activeMask = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  perLaneConflictReq_reg_7_bankIdx = _RAND_17[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_11(
  input        clock,
  input        reset,
  input        io_r_req_valid,
  input  [6:0] io_r_req_bits_setIdx,
  output [7:0] io_r_resp_data_0,
  output [7:0] io_r_resp_data_1,
  output [7:0] io_r_resp_data_2,
  output [7:0] io_r_resp_data_3,
  input        io_w_req_valid,
  input  [6:0] io_w_req_bits_setIdx,
  input  [7:0] io_w_req_bits_data_0,
  input  [7:0] io_w_req_bits_data_1,
  input  [7:0] io_w_req_bits_data_2,
  input  [7:0] io_w_req_bits_data_3,
  input  [3:0] io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] array_0 [0:127]; // @[SRAMTemplate.scala 101:26]
  wire  array_0_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_0_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_0_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_0_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_0_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_0_raw_rdata_en_pipe_0;
  reg [6:0] array_0_raw_rdata_addr_pipe_0;
  reg [7:0] array_1 [0:127]; // @[SRAMTemplate.scala 101:26]
  wire  array_1_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_1_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_1_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_1_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_1_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_1_raw_rdata_en_pipe_0;
  reg [6:0] array_1_raw_rdata_addr_pipe_0;
  reg [7:0] array_2 [0:127]; // @[SRAMTemplate.scala 101:26]
  wire  array_2_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_2_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_2_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_2_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_2_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_2_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_2_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_2_raw_rdata_en_pipe_0;
  reg [6:0] array_2_raw_rdata_addr_pipe_0;
  reg [7:0] array_3 [0:127]; // @[SRAMTemplate.scala 101:26]
  wire  array_3_raw_rdata_en; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_3_raw_rdata_addr; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_3_raw_rdata_data; // @[SRAMTemplate.scala 101:26]
  wire [7:0] array_3_MPORT_data; // @[SRAMTemplate.scala 101:26]
  wire [6:0] array_3_MPORT_addr; // @[SRAMTemplate.scala 101:26]
  wire  array_3_MPORT_mask; // @[SRAMTemplate.scala 101:26]
  wire  array_3_MPORT_en; // @[SRAMTemplate.scala 101:26]
  reg  array_3_raw_rdata_en_pipe_0;
  reg [6:0] array_3_raw_rdata_addr_pipe_0;
  reg [63:0] bypass_wdata_lfsr; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor = bypass_wdata_lfsr[0] ^ bypass_wdata_lfsr[1] ^ bypass_wdata_lfsr[3] ^ bypass_wdata_lfsr[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_2 = {bypass_wdata_xor,bypass_wdata_lfsr[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_1; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_1 = bypass_wdata_lfsr_1[0] ^ bypass_wdata_lfsr_1[1] ^ bypass_wdata_lfsr_1[3] ^
    bypass_wdata_lfsr_1[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_6 = {bypass_wdata_xor_1,bypass_wdata_lfsr_1[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_2; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_2 = bypass_wdata_lfsr_2[0] ^ bypass_wdata_lfsr_2[1] ^ bypass_wdata_lfsr_2[3] ^
    bypass_wdata_lfsr_2[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_10 = {bypass_wdata_xor_2,bypass_wdata_lfsr_2[63:1]}; // @[Cat.scala 31:58]
  reg [63:0] bypass_wdata_lfsr_3; // @[LFSR64.scala 25:23]
  wire  bypass_wdata_xor_3 = bypass_wdata_lfsr_3[0] ^ bypass_wdata_lfsr_3[1] ^ bypass_wdata_lfsr_3[3] ^
    bypass_wdata_lfsr_3[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _bypass_wdata_lfsr_T_14 = {bypass_wdata_xor_3,bypass_wdata_lfsr_3[63:1]}; // @[Cat.scala 31:58]
  reg  bypass_mask_need_check; // @[SRAMTemplate.scala 126:29]
  reg [6:0] bypass_mask_waddr_reg; // @[SRAMTemplate.scala 127:28]
  reg [6:0] bypass_mask_raddr_reg; // @[SRAMTemplate.scala 128:28]
  wire  _bypass_mask_bypass_T_1 = bypass_mask_need_check & bypass_mask_waddr_reg == bypass_mask_raddr_reg; // @[SRAMTemplate.scala 130:39]
  wire [3:0] _bypass_mask_bypass_T_3 = _bypass_mask_bypass_T_1 ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  reg [3:0] bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:76]
  wire [3:0] bypass_mask_bypass = _bypass_mask_bypass_T_3 & bypass_mask_bypass_REG; // @[SRAMTemplate.scala 130:67]
  wire [7:0] bypass_wdata_0 = bypass_wdata_lfsr[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [7:0] bypass_wdata_1 = bypass_wdata_lfsr_1[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [7:0] bypass_wdata_2 = bypass_wdata_lfsr_2[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  wire [7:0] bypass_wdata_3 = bypass_wdata_lfsr_3[7:0]; // @[SRAMTemplate.scala 134:{58,58}]
  assign array_0_raw_rdata_en = array_0_raw_rdata_en_pipe_0;
  assign array_0_raw_rdata_addr = array_0_raw_rdata_addr_pipe_0;
  assign array_0_raw_rdata_data = array_0[array_0_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_0_MPORT_data = io_w_req_bits_data_0;
  assign array_0_MPORT_addr = io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = io_w_req_bits_waymask[0];
  assign array_0_MPORT_en = io_w_req_valid;
  assign array_1_raw_rdata_en = array_1_raw_rdata_en_pipe_0;
  assign array_1_raw_rdata_addr = array_1_raw_rdata_addr_pipe_0;
  assign array_1_raw_rdata_data = array_1[array_1_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_1_MPORT_data = io_w_req_bits_data_1;
  assign array_1_MPORT_addr = io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = io_w_req_bits_waymask[1];
  assign array_1_MPORT_en = io_w_req_valid;
  assign array_2_raw_rdata_en = array_2_raw_rdata_en_pipe_0;
  assign array_2_raw_rdata_addr = array_2_raw_rdata_addr_pipe_0;
  assign array_2_raw_rdata_data = array_2[array_2_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_2_MPORT_data = io_w_req_bits_data_2;
  assign array_2_MPORT_addr = io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = io_w_req_bits_waymask[2];
  assign array_2_MPORT_en = io_w_req_valid;
  assign array_3_raw_rdata_en = array_3_raw_rdata_en_pipe_0;
  assign array_3_raw_rdata_addr = array_3_raw_rdata_addr_pipe_0;
  assign array_3_raw_rdata_data = array_3[array_3_raw_rdata_addr]; // @[SRAMTemplate.scala 101:26]
  assign array_3_MPORT_data = io_w_req_bits_data_3;
  assign array_3_MPORT_addr = io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = io_w_req_bits_waymask[3];
  assign array_3_MPORT_en = io_w_req_valid;
  assign io_r_resp_data_0 = bypass_mask_bypass[0] ? bypass_wdata_0 : array_0_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_1 = bypass_mask_bypass[1] ? bypass_wdata_1 : array_1_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_2 = bypass_mask_bypass[2] ? bypass_wdata_2 : array_2_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  assign io_r_resp_data_3 = bypass_mask_bypass[3] ? bypass_wdata_3 : array_3_raw_rdata_data; // @[SRAMTemplate.scala 139:30]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_0_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_0_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_1_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_1_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_2_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_2_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[SRAMTemplate.scala 101:26]
    end
    array_3_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_3_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr <= 64'h1;
    end else begin
      bypass_wdata_lfsr <= _bypass_wdata_lfsr_T_2;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_1 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_1 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_1 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_1 <= _bypass_wdata_lfsr_T_6;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_2 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_2 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_2 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_2 <= _bypass_wdata_lfsr_T_10;
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      bypass_wdata_lfsr_3 <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (bypass_wdata_lfsr_3 == 64'h0) begin // @[LFSR64.scala 28:18]
      bypass_wdata_lfsr_3 <= 64'h1;
    end else begin
      bypass_wdata_lfsr_3 <= _bypass_wdata_lfsr_T_14;
    end
    bypass_mask_need_check <= io_r_req_valid & io_w_req_valid; // @[SRAMTemplate.scala 126:34]
    bypass_mask_waddr_reg <= io_w_req_bits_setIdx; // @[SRAMTemplate.scala 127:28]
    bypass_mask_raddr_reg <= io_r_req_bits_setIdx; // @[SRAMTemplate.scala 128:28]
    bypass_mask_bypass_REG <= io_w_req_bits_waymask; // @[SRAMTemplate.scala 130:76]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_3[initvar] = _RAND_9[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_raw_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_raw_rdata_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_raw_rdata_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_raw_rdata_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_raw_rdata_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_raw_rdata_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_raw_rdata_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_raw_rdata_addr_pipe_0 = _RAND_11[6:0];
  _RAND_12 = {2{`RANDOM}};
  bypass_wdata_lfsr = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  bypass_wdata_lfsr_1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  bypass_wdata_lfsr_2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  bypass_wdata_lfsr_3 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  bypass_mask_need_check = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  bypass_mask_waddr_reg = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  bypass_mask_raddr_reg = _RAND_18[6:0];
  _RAND_19 = {1{`RANDOM}};
  bypass_mask_bypass_REG = _RAND_19[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SharedMemory(
  input         clock,
  input         reset,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [1:0]  io_coreReq_bits_instrId,
  input         io_coreReq_bits_isWrite,
  input  [6:0]  io_coreReq_bits_setIdx,
  input         io_coreReq_bits_perLaneAddr_0_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_0_blockOffset,
  input         io_coreReq_bits_perLaneAddr_1_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_1_blockOffset,
  input         io_coreReq_bits_perLaneAddr_2_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_2_blockOffset,
  input         io_coreReq_bits_perLaneAddr_3_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_3_blockOffset,
  input         io_coreReq_bits_perLaneAddr_4_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_4_blockOffset,
  input         io_coreReq_bits_perLaneAddr_5_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_5_blockOffset,
  input         io_coreReq_bits_perLaneAddr_6_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_6_blockOffset,
  input         io_coreReq_bits_perLaneAddr_7_activeMask,
  input  [2:0]  io_coreReq_bits_perLaneAddr_7_blockOffset,
  input  [31:0] io_coreReq_bits_data_0,
  input  [31:0] io_coreReq_bits_data_1,
  input  [31:0] io_coreReq_bits_data_2,
  input  [31:0] io_coreReq_bits_data_3,
  input  [31:0] io_coreReq_bits_data_4,
  input  [31:0] io_coreReq_bits_data_5,
  input  [31:0] io_coreReq_bits_data_6,
  input  [31:0] io_coreReq_bits_data_7,
  input         io_coreRsp_ready,
  output        io_coreRsp_valid,
  output [1:0]  io_coreRsp_bits_instrId,
  output [31:0] io_coreRsp_bits_data_0,
  output [31:0] io_coreRsp_bits_data_1,
  output [31:0] io_coreRsp_bits_data_2,
  output [31:0] io_coreRsp_bits_data_3,
  output [31:0] io_coreRsp_bits_data_4,
  output [31:0] io_coreRsp_bits_data_5,
  output [31:0] io_coreRsp_bits_data_6,
  output [31:0] io_coreRsp_bits_data_7,
  output        io_coreRsp_bits_activeMask_0,
  output        io_coreRsp_bits_activeMask_1,
  output        io_coreRsp_bits_activeMask_2,
  output        io_coreRsp_bits_activeMask_3,
  output        io_coreRsp_bits_activeMask_4,
  output        io_coreRsp_bits_activeMask_5,
  output        io_coreRsp_bits_activeMask_6,
  output        io_coreRsp_bits_activeMask_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
`endif // RANDOMIZE_REG_INIT
  wire  BankConfArb_clock; // @[ShareMem.scala 46:27]
  wire  BankConfArb_reset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_isWrite; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_0_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_0_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_1_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_1_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_2_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_2_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_3_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_3_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_4_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_4_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_5_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_5_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_6_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_6_blockOffset; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_coreReqArb_perLaneAddr_7_activeMask; // @[ShareMem.scala 46:27]
  wire [2:0] BankConfArb_io_coreReqArb_perLaneAddr_7_blockOffset; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_0; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_1; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_2; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_3; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_4; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_5; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_6; // @[ShareMem.scala 46:27]
  wire [7:0] BankConfArb_io_dataCrsbarSel1H_7; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_0_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_1_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_2_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_3_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_4_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_5_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_6_wordOffset1H; // @[ShareMem.scala 46:27]
  wire [3:0] BankConfArb_io_addrCrsbarOut_7_wordOffset1H; // @[ShareMem.scala 46:27]
  wire  BankConfArb_io_bankConflict; // @[ShareMem.scala 46:27]
  wire [31:0] DataCorssBarForWrite_io_DataIn_0; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_1; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_2; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_3; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_4; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_5; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_6; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataIn_7; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_0; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_1; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_2; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_3; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_4; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_5; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_6; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForWrite_io_DataOut_7; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_0; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_1; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_2; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_3; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_4; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_5; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_6; // @[ShareMem.scala 48:36]
  wire [7:0] DataCorssBarForWrite_io_Select1H_7; // @[ShareMem.scala 48:36]
  wire [31:0] DataCorssBarForRead_io_DataIn_0; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_1; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_2; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_3; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_4; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_5; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_6; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataIn_7; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_0; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_1; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_2; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_3; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_4; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_5; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_6; // @[ShareMem.scala 49:35]
  wire [31:0] DataCorssBarForRead_io_DataOut_7; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_0; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_1; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_2; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_3; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_4; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_5; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_6; // @[ShareMem.scala 49:35]
  wire [7:0] DataCorssBarForRead_io_Select1H_7; // @[ShareMem.scala 49:35]
  wire  coreRsp_Q_clock; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_reset; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_ready; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_valid; // @[ShareMem.scala 57:25]
  wire [1:0] coreRsp_Q_io_enq_bits_instrId; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_0; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_1; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_2; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_3; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_4; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_5; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_6; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_enq_bits_data_7; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_0; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_1; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_2; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_3; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_4; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_5; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_6; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_enq_bits_activeMask_7; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_ready; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_valid; // @[ShareMem.scala 57:25]
  wire [1:0] coreRsp_Q_io_deq_bits_instrId; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_0; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_1; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_2; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_3; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_4; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_5; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_6; // @[ShareMem.scala 57:25]
  wire [31:0] coreRsp_Q_io_deq_bits_data_7; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_0; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_1; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_2; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_3; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_4; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_5; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_6; // @[ShareMem.scala 57:25]
  wire  coreRsp_Q_io_deq_bits_activeMask_7; // @[ShareMem.scala 57:25]
  wire [2:0] coreRsp_Q_io_count; // @[ShareMem.scala 57:25]
  wire  DataAccessesRRsp_DataAccess_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_1_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_1_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_1_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_1_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_1_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_1_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_2_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_2_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_2_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_2_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_2_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_2_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_3_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_3_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_3_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_3_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_3_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_3_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_4_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_4_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_4_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_4_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_4_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_4_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_5_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_5_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_5_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_5_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_5_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_5_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_6_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_6_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_6_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_6_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_6_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_6_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_7_clock; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_7_reset; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_7_io_r_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_7_io_r_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_r_resp_data_3; // @[ShareMem.scala 123:28]
  wire  DataAccessesRRsp_DataAccess_7_io_w_req_valid; // @[ShareMem.scala 123:28]
  wire [6:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_setIdx; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_0; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_1; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_2; // @[ShareMem.scala 123:28]
  wire [7:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_3; // @[ShareMem.scala 123:28]
  wire [3:0] DataAccessesRRsp_DataAccess_7_io_w_req_bits_waymask; // @[ShareMem.scala 123:28]
  wire  _coreReqisValidWrite_st1_T = io_coreReq_ready & io_coreReq_valid; // @[Decoupled.scala 50:35]
  reg  coreReqisValidWrite_st1; // @[ShareMem.scala 103:40]
  wire  _coreReqisValidRead_st1_T_1 = ~io_coreReq_bits_isWrite; // @[ShareMem.scala 104:62]
  reg  coreReqisValidRead_st1; // @[ShareMem.scala 104:40]
  reg  coreReqisValidRead_st2; // @[ShareMem.scala 105:39]
  reg  coreReqisValidWrite_st2; // @[ShareMem.scala 106:40]
  reg [1:0] coreReq_st1_instrId; // @[Reg.scala 16:16]
  reg [6:0] coreReq_st1_setIdx; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_0_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_1_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_2_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_3_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_4_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_5_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_6_activeMask; // @[Reg.scala 16:16]
  reg  coreReq_st1_perLaneAddr_7_activeMask; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_0; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_1; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_2; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_3; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_4; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_5; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_6; // @[Reg.scala 16:16]
  reg [31:0] coreReq_st1_data_7; // @[Reg.scala 16:16]
  reg [1:0] coreReqInstrId_st2; // @[ShareMem.scala 109:35]
  reg  coreReqActvMask_st2_0; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_1; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_2; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_3; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_4; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_5; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_6; // @[ShareMem.scala 110:36]
  reg  coreReqActvMask_st2_7; // @[ShareMem.scala 110:36]
  reg [3:0] arbAddrCrsbarOut_st1_0_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_1_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_2_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_3_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_4_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_5_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_6_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [3:0] arbAddrCrsbarOut_st1_7_wordOffset1H; // @[ShareMem.scala 113:37]
  reg [7:0] arbDataCrsbarSel1H_st1_0; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_1; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_2; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_3; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_4; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_5; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_6; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st1_7; // @[ShareMem.scala 114:39]
  reg [7:0] arbDataCrsbarSel1H_st2_0; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_1; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_2; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_3; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_4; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_5; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_6; // @[ShareMem.scala 115:39]
  reg [7:0] arbDataCrsbarSel1H_st2_7; // @[ShareMem.scala 115:39]
  wire [31:0] _DataAccessesRRsp_WIRE_1 = DataCorssBarForWrite_io_DataOut_0;
  wire [31:0] DataAccessesRRsp_0 = {DataAccessesRRsp_DataAccess_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_io_r_resp_data_2,DataAccessesRRsp_DataAccess_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_3 = DataCorssBarForWrite_io_DataOut_1;
  wire [31:0] DataAccessesRRsp_1 = {DataAccessesRRsp_DataAccess_1_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_1_io_r_resp_data_2,DataAccessesRRsp_DataAccess_1_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_1_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_5 = DataCorssBarForWrite_io_DataOut_2;
  wire [31:0] DataAccessesRRsp_2 = {DataAccessesRRsp_DataAccess_2_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_2_io_r_resp_data_2,DataAccessesRRsp_DataAccess_2_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_2_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_7 = DataCorssBarForWrite_io_DataOut_3;
  wire [31:0] DataAccessesRRsp_3 = {DataAccessesRRsp_DataAccess_3_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_3_io_r_resp_data_2,DataAccessesRRsp_DataAccess_3_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_3_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_9 = DataCorssBarForWrite_io_DataOut_4;
  wire [31:0] DataAccessesRRsp_4 = {DataAccessesRRsp_DataAccess_4_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_4_io_r_resp_data_2,DataAccessesRRsp_DataAccess_4_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_4_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_11 = DataCorssBarForWrite_io_DataOut_5;
  wire [31:0] DataAccessesRRsp_5 = {DataAccessesRRsp_DataAccess_5_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_5_io_r_resp_data_2,DataAccessesRRsp_DataAccess_5_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_5_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_13 = DataCorssBarForWrite_io_DataOut_6;
  wire [31:0] DataAccessesRRsp_6 = {DataAccessesRRsp_DataAccess_6_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_6_io_r_resp_data_2,DataAccessesRRsp_DataAccess_6_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_6_io_r_resp_data_0}; // @[Cat.scala 31:58]
  wire [31:0] _DataAccessesRRsp_WIRE_15 = DataCorssBarForWrite_io_DataOut_7;
  wire [31:0] DataAccessesRRsp_7 = {DataAccessesRRsp_DataAccess_7_io_r_resp_data_3,
    DataAccessesRRsp_DataAccess_7_io_r_resp_data_2,DataAccessesRRsp_DataAccess_7_io_r_resp_data_1,
    DataAccessesRRsp_DataAccess_7_io_r_resp_data_0}; // @[Cat.scala 31:58]
  reg [31:0] dataAccess_data_st2_0; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_1; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_2; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_3; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_4; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_5; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_6; // @[Reg.scala 16:16]
  reg [31:0] dataAccess_data_st2_7; // @[Reg.scala 16:16]
  wire [2:0] _coreRsp_QAlmstFull_T_1 = 3'h4 - 3'h2; // @[ShareMem.scala 166:70]
  wire  coreRsp_QAlmstFull = coreRsp_Q_io_count == _coreRsp_QAlmstFull_T_1; // @[ShareMem.scala 166:44]
  BankConflictArbiter_1 BankConfArb ( // @[ShareMem.scala 46:27]
    .clock(BankConfArb_clock),
    .reset(BankConfArb_reset),
    .io_coreReqArb_isWrite(BankConfArb_io_coreReqArb_isWrite),
    .io_coreReqArb_perLaneAddr_0_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_0_activeMask),
    .io_coreReqArb_perLaneAddr_0_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_0_blockOffset),
    .io_coreReqArb_perLaneAddr_1_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_1_activeMask),
    .io_coreReqArb_perLaneAddr_1_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_1_blockOffset),
    .io_coreReqArb_perLaneAddr_2_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_2_activeMask),
    .io_coreReqArb_perLaneAddr_2_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_2_blockOffset),
    .io_coreReqArb_perLaneAddr_3_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_3_activeMask),
    .io_coreReqArb_perLaneAddr_3_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_3_blockOffset),
    .io_coreReqArb_perLaneAddr_4_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_4_activeMask),
    .io_coreReqArb_perLaneAddr_4_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_4_blockOffset),
    .io_coreReqArb_perLaneAddr_5_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_5_activeMask),
    .io_coreReqArb_perLaneAddr_5_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_5_blockOffset),
    .io_coreReqArb_perLaneAddr_6_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_6_activeMask),
    .io_coreReqArb_perLaneAddr_6_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_6_blockOffset),
    .io_coreReqArb_perLaneAddr_7_activeMask(BankConfArb_io_coreReqArb_perLaneAddr_7_activeMask),
    .io_coreReqArb_perLaneAddr_7_blockOffset(BankConfArb_io_coreReqArb_perLaneAddr_7_blockOffset),
    .io_dataCrsbarSel1H_0(BankConfArb_io_dataCrsbarSel1H_0),
    .io_dataCrsbarSel1H_1(BankConfArb_io_dataCrsbarSel1H_1),
    .io_dataCrsbarSel1H_2(BankConfArb_io_dataCrsbarSel1H_2),
    .io_dataCrsbarSel1H_3(BankConfArb_io_dataCrsbarSel1H_3),
    .io_dataCrsbarSel1H_4(BankConfArb_io_dataCrsbarSel1H_4),
    .io_dataCrsbarSel1H_5(BankConfArb_io_dataCrsbarSel1H_5),
    .io_dataCrsbarSel1H_6(BankConfArb_io_dataCrsbarSel1H_6),
    .io_dataCrsbarSel1H_7(BankConfArb_io_dataCrsbarSel1H_7),
    .io_addrCrsbarOut_0_wordOffset1H(BankConfArb_io_addrCrsbarOut_0_wordOffset1H),
    .io_addrCrsbarOut_1_wordOffset1H(BankConfArb_io_addrCrsbarOut_1_wordOffset1H),
    .io_addrCrsbarOut_2_wordOffset1H(BankConfArb_io_addrCrsbarOut_2_wordOffset1H),
    .io_addrCrsbarOut_3_wordOffset1H(BankConfArb_io_addrCrsbarOut_3_wordOffset1H),
    .io_addrCrsbarOut_4_wordOffset1H(BankConfArb_io_addrCrsbarOut_4_wordOffset1H),
    .io_addrCrsbarOut_5_wordOffset1H(BankConfArb_io_addrCrsbarOut_5_wordOffset1H),
    .io_addrCrsbarOut_6_wordOffset1H(BankConfArb_io_addrCrsbarOut_6_wordOffset1H),
    .io_addrCrsbarOut_7_wordOffset1H(BankConfArb_io_addrCrsbarOut_7_wordOffset1H),
    .io_bankConflict(BankConfArb_io_bankConflict)
  );
  DataCrossbar DataCorssBarForWrite ( // @[ShareMem.scala 48:36]
    .io_DataIn_0(DataCorssBarForWrite_io_DataIn_0),
    .io_DataIn_1(DataCorssBarForWrite_io_DataIn_1),
    .io_DataIn_2(DataCorssBarForWrite_io_DataIn_2),
    .io_DataIn_3(DataCorssBarForWrite_io_DataIn_3),
    .io_DataIn_4(DataCorssBarForWrite_io_DataIn_4),
    .io_DataIn_5(DataCorssBarForWrite_io_DataIn_5),
    .io_DataIn_6(DataCorssBarForWrite_io_DataIn_6),
    .io_DataIn_7(DataCorssBarForWrite_io_DataIn_7),
    .io_DataOut_0(DataCorssBarForWrite_io_DataOut_0),
    .io_DataOut_1(DataCorssBarForWrite_io_DataOut_1),
    .io_DataOut_2(DataCorssBarForWrite_io_DataOut_2),
    .io_DataOut_3(DataCorssBarForWrite_io_DataOut_3),
    .io_DataOut_4(DataCorssBarForWrite_io_DataOut_4),
    .io_DataOut_5(DataCorssBarForWrite_io_DataOut_5),
    .io_DataOut_6(DataCorssBarForWrite_io_DataOut_6),
    .io_DataOut_7(DataCorssBarForWrite_io_DataOut_7),
    .io_Select1H_0(DataCorssBarForWrite_io_Select1H_0),
    .io_Select1H_1(DataCorssBarForWrite_io_Select1H_1),
    .io_Select1H_2(DataCorssBarForWrite_io_Select1H_2),
    .io_Select1H_3(DataCorssBarForWrite_io_Select1H_3),
    .io_Select1H_4(DataCorssBarForWrite_io_Select1H_4),
    .io_Select1H_5(DataCorssBarForWrite_io_Select1H_5),
    .io_Select1H_6(DataCorssBarForWrite_io_Select1H_6),
    .io_Select1H_7(DataCorssBarForWrite_io_Select1H_7)
  );
  DataCrossbar DataCorssBarForRead ( // @[ShareMem.scala 49:35]
    .io_DataIn_0(DataCorssBarForRead_io_DataIn_0),
    .io_DataIn_1(DataCorssBarForRead_io_DataIn_1),
    .io_DataIn_2(DataCorssBarForRead_io_DataIn_2),
    .io_DataIn_3(DataCorssBarForRead_io_DataIn_3),
    .io_DataIn_4(DataCorssBarForRead_io_DataIn_4),
    .io_DataIn_5(DataCorssBarForRead_io_DataIn_5),
    .io_DataIn_6(DataCorssBarForRead_io_DataIn_6),
    .io_DataIn_7(DataCorssBarForRead_io_DataIn_7),
    .io_DataOut_0(DataCorssBarForRead_io_DataOut_0),
    .io_DataOut_1(DataCorssBarForRead_io_DataOut_1),
    .io_DataOut_2(DataCorssBarForRead_io_DataOut_2),
    .io_DataOut_3(DataCorssBarForRead_io_DataOut_3),
    .io_DataOut_4(DataCorssBarForRead_io_DataOut_4),
    .io_DataOut_5(DataCorssBarForRead_io_DataOut_5),
    .io_DataOut_6(DataCorssBarForRead_io_DataOut_6),
    .io_DataOut_7(DataCorssBarForRead_io_DataOut_7),
    .io_Select1H_0(DataCorssBarForRead_io_Select1H_0),
    .io_Select1H_1(DataCorssBarForRead_io_Select1H_1),
    .io_Select1H_2(DataCorssBarForRead_io_Select1H_2),
    .io_Select1H_3(DataCorssBarForRead_io_Select1H_3),
    .io_Select1H_4(DataCorssBarForRead_io_Select1H_4),
    .io_Select1H_5(DataCorssBarForRead_io_Select1H_5),
    .io_Select1H_6(DataCorssBarForRead_io_Select1H_6),
    .io_Select1H_7(DataCorssBarForRead_io_Select1H_7)
  );
  Queue_50 coreRsp_Q ( // @[ShareMem.scala 57:25]
    .clock(coreRsp_Q_clock),
    .reset(coreRsp_Q_reset),
    .io_enq_ready(coreRsp_Q_io_enq_ready),
    .io_enq_valid(coreRsp_Q_io_enq_valid),
    .io_enq_bits_instrId(coreRsp_Q_io_enq_bits_instrId),
    .io_enq_bits_data_0(coreRsp_Q_io_enq_bits_data_0),
    .io_enq_bits_data_1(coreRsp_Q_io_enq_bits_data_1),
    .io_enq_bits_data_2(coreRsp_Q_io_enq_bits_data_2),
    .io_enq_bits_data_3(coreRsp_Q_io_enq_bits_data_3),
    .io_enq_bits_data_4(coreRsp_Q_io_enq_bits_data_4),
    .io_enq_bits_data_5(coreRsp_Q_io_enq_bits_data_5),
    .io_enq_bits_data_6(coreRsp_Q_io_enq_bits_data_6),
    .io_enq_bits_data_7(coreRsp_Q_io_enq_bits_data_7),
    .io_enq_bits_activeMask_0(coreRsp_Q_io_enq_bits_activeMask_0),
    .io_enq_bits_activeMask_1(coreRsp_Q_io_enq_bits_activeMask_1),
    .io_enq_bits_activeMask_2(coreRsp_Q_io_enq_bits_activeMask_2),
    .io_enq_bits_activeMask_3(coreRsp_Q_io_enq_bits_activeMask_3),
    .io_enq_bits_activeMask_4(coreRsp_Q_io_enq_bits_activeMask_4),
    .io_enq_bits_activeMask_5(coreRsp_Q_io_enq_bits_activeMask_5),
    .io_enq_bits_activeMask_6(coreRsp_Q_io_enq_bits_activeMask_6),
    .io_enq_bits_activeMask_7(coreRsp_Q_io_enq_bits_activeMask_7),
    .io_deq_ready(coreRsp_Q_io_deq_ready),
    .io_deq_valid(coreRsp_Q_io_deq_valid),
    .io_deq_bits_instrId(coreRsp_Q_io_deq_bits_instrId),
    .io_deq_bits_data_0(coreRsp_Q_io_deq_bits_data_0),
    .io_deq_bits_data_1(coreRsp_Q_io_deq_bits_data_1),
    .io_deq_bits_data_2(coreRsp_Q_io_deq_bits_data_2),
    .io_deq_bits_data_3(coreRsp_Q_io_deq_bits_data_3),
    .io_deq_bits_data_4(coreRsp_Q_io_deq_bits_data_4),
    .io_deq_bits_data_5(coreRsp_Q_io_deq_bits_data_5),
    .io_deq_bits_data_6(coreRsp_Q_io_deq_bits_data_6),
    .io_deq_bits_data_7(coreRsp_Q_io_deq_bits_data_7),
    .io_deq_bits_activeMask_0(coreRsp_Q_io_deq_bits_activeMask_0),
    .io_deq_bits_activeMask_1(coreRsp_Q_io_deq_bits_activeMask_1),
    .io_deq_bits_activeMask_2(coreRsp_Q_io_deq_bits_activeMask_2),
    .io_deq_bits_activeMask_3(coreRsp_Q_io_deq_bits_activeMask_3),
    .io_deq_bits_activeMask_4(coreRsp_Q_io_deq_bits_activeMask_4),
    .io_deq_bits_activeMask_5(coreRsp_Q_io_deq_bits_activeMask_5),
    .io_deq_bits_activeMask_6(coreRsp_Q_io_deq_bits_activeMask_6),
    .io_deq_bits_activeMask_7(coreRsp_Q_io_deq_bits_activeMask_7),
    .io_count(coreRsp_Q_io_count)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_clock),
    .reset(DataAccessesRRsp_DataAccess_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_1 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_1_clock),
    .reset(DataAccessesRRsp_DataAccess_1_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_1_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_1_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_1_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_1_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_1_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_1_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_1_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_1_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_1_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_2 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_2_clock),
    .reset(DataAccessesRRsp_DataAccess_2_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_2_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_2_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_2_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_2_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_2_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_2_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_2_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_2_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_2_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_3 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_3_clock),
    .reset(DataAccessesRRsp_DataAccess_3_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_3_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_3_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_3_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_3_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_3_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_3_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_3_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_3_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_3_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_4 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_4_clock),
    .reset(DataAccessesRRsp_DataAccess_4_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_4_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_4_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_4_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_4_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_4_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_4_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_4_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_4_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_4_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_5 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_5_clock),
    .reset(DataAccessesRRsp_DataAccess_5_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_5_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_5_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_5_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_5_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_5_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_5_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_5_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_5_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_5_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_6 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_6_clock),
    .reset(DataAccessesRRsp_DataAccess_6_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_6_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_6_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_6_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_6_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_6_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_6_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_6_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_6_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_6_io_w_req_bits_waymask)
  );
  SRAMTemplate_11 DataAccessesRRsp_DataAccess_7 ( // @[ShareMem.scala 123:28]
    .clock(DataAccessesRRsp_DataAccess_7_clock),
    .reset(DataAccessesRRsp_DataAccess_7_reset),
    .io_r_req_valid(DataAccessesRRsp_DataAccess_7_io_r_req_valid),
    .io_r_req_bits_setIdx(DataAccessesRRsp_DataAccess_7_io_r_req_bits_setIdx),
    .io_r_resp_data_0(DataAccessesRRsp_DataAccess_7_io_r_resp_data_0),
    .io_r_resp_data_1(DataAccessesRRsp_DataAccess_7_io_r_resp_data_1),
    .io_r_resp_data_2(DataAccessesRRsp_DataAccess_7_io_r_resp_data_2),
    .io_r_resp_data_3(DataAccessesRRsp_DataAccess_7_io_r_resp_data_3),
    .io_w_req_valid(DataAccessesRRsp_DataAccess_7_io_w_req_valid),
    .io_w_req_bits_setIdx(DataAccessesRRsp_DataAccess_7_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(DataAccessesRRsp_DataAccess_7_io_w_req_bits_waymask)
  );
  assign io_coreReq_ready = ~BankConfArb_io_bankConflict & ~coreRsp_QAlmstFull; // @[ShareMem.scala 170:52]
  assign io_coreRsp_valid = coreRsp_Q_io_deq_valid; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_instrId = coreRsp_Q_io_deq_bits_instrId; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_0 = coreRsp_Q_io_deq_bits_data_0; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_1 = coreRsp_Q_io_deq_bits_data_1; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_2 = coreRsp_Q_io_deq_bits_data_2; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_3 = coreRsp_Q_io_deq_bits_data_3; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_4 = coreRsp_Q_io_deq_bits_data_4; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_5 = coreRsp_Q_io_deq_bits_data_5; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_6 = coreRsp_Q_io_deq_bits_data_6; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_data_7 = coreRsp_Q_io_deq_bits_data_7; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_0 = coreRsp_Q_io_deq_bits_activeMask_0; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_1 = coreRsp_Q_io_deq_bits_activeMask_1; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_2 = coreRsp_Q_io_deq_bits_activeMask_2; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_3 = coreRsp_Q_io_deq_bits_activeMask_3; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_4 = coreRsp_Q_io_deq_bits_activeMask_4; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_5 = coreRsp_Q_io_deq_bits_activeMask_5; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_6 = coreRsp_Q_io_deq_bits_activeMask_6; // @[ShareMem.scala 160:20]
  assign io_coreRsp_bits_activeMask_7 = coreRsp_Q_io_deq_bits_activeMask_7; // @[ShareMem.scala 160:20]
  assign BankConfArb_clock = clock;
  assign BankConfArb_reset = reset;
  assign BankConfArb_io_coreReqArb_isWrite = io_coreReq_bits_isWrite; // @[ShareMem.scala 62:37]
  assign BankConfArb_io_coreReqArb_perLaneAddr_0_activeMask = io_coreReq_bits_perLaneAddr_0_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_0_blockOffset = io_coreReq_bits_perLaneAddr_0_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_1_activeMask = io_coreReq_bits_perLaneAddr_1_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_1_blockOffset = io_coreReq_bits_perLaneAddr_1_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_2_activeMask = io_coreReq_bits_perLaneAddr_2_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_2_blockOffset = io_coreReq_bits_perLaneAddr_2_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_3_activeMask = io_coreReq_bits_perLaneAddr_3_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_3_blockOffset = io_coreReq_bits_perLaneAddr_3_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_4_activeMask = io_coreReq_bits_perLaneAddr_4_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_4_blockOffset = io_coreReq_bits_perLaneAddr_4_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_5_activeMask = io_coreReq_bits_perLaneAddr_5_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_5_blockOffset = io_coreReq_bits_perLaneAddr_5_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_6_activeMask = io_coreReq_bits_perLaneAddr_6_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_6_blockOffset = io_coreReq_bits_perLaneAddr_6_blockOffset; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_7_activeMask = io_coreReq_bits_perLaneAddr_7_activeMask; // @[ShareMem.scala 63:41]
  assign BankConfArb_io_coreReqArb_perLaneAddr_7_blockOffset = io_coreReq_bits_perLaneAddr_7_blockOffset; // @[ShareMem.scala 63:41]
  assign DataCorssBarForWrite_io_DataIn_0 = coreReq_st1_data_0; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_1 = coreReq_st1_data_1; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_2 = coreReq_st1_data_2; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_3 = coreReq_st1_data_3; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_4 = coreReq_st1_data_4; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_5 = coreReq_st1_data_5; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_6 = coreReq_st1_data_6; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_DataIn_7 = coreReq_st1_data_7; // @[ShareMem.scala 153:34]
  assign DataCorssBarForWrite_io_Select1H_0 = arbDataCrsbarSel1H_st1_0; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_1 = arbDataCrsbarSel1H_st1_1; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_2 = arbDataCrsbarSel1H_st1_2; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_3 = arbDataCrsbarSel1H_st1_3; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_4 = arbDataCrsbarSel1H_st1_4; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_5 = arbDataCrsbarSel1H_st1_5; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_6 = arbDataCrsbarSel1H_st1_6; // @[ShareMem.scala 154:36]
  assign DataCorssBarForWrite_io_Select1H_7 = arbDataCrsbarSel1H_st1_7; // @[ShareMem.scala 154:36]
  assign DataCorssBarForRead_io_DataIn_0 = dataAccess_data_st2_0; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_1 = dataAccess_data_st2_1; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_2 = dataAccess_data_st2_2; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_3 = dataAccess_data_st2_3; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_4 = dataAccess_data_st2_4; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_5 = dataAccess_data_st2_5; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_6 = dataAccess_data_st2_6; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_DataIn_7 = dataAccess_data_st2_7; // @[ShareMem.scala 156:33]
  assign DataCorssBarForRead_io_Select1H_0 = arbDataCrsbarSel1H_st2_0; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_1 = arbDataCrsbarSel1H_st2_1; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_2 = arbDataCrsbarSel1H_st2_2; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_3 = arbDataCrsbarSel1H_st2_3; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_4 = arbDataCrsbarSel1H_st2_4; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_5 = arbDataCrsbarSel1H_st2_5; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_6 = arbDataCrsbarSel1H_st2_6; // @[ShareMem.scala 157:35]
  assign DataCorssBarForRead_io_Select1H_7 = arbDataCrsbarSel1H_st2_7; // @[ShareMem.scala 157:35]
  assign coreRsp_Q_clock = clock;
  assign coreRsp_Q_reset = reset;
  assign coreRsp_Q_io_enq_valid = coreReqisValidRead_st2 | coreReqisValidWrite_st2; // @[ShareMem.scala 161:52]
  assign coreRsp_Q_io_enq_bits_instrId = coreReqInstrId_st2; // @[ShareMem.scala 164:33]
  assign coreRsp_Q_io_enq_bits_data_0 = DataCorssBarForRead_io_DataOut_0; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_1 = DataCorssBarForRead_io_DataOut_1; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_2 = DataCorssBarForRead_io_DataOut_2; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_3 = DataCorssBarForRead_io_DataOut_3; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_4 = DataCorssBarForRead_io_DataOut_4; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_5 = DataCorssBarForRead_io_DataOut_5; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_6 = DataCorssBarForRead_io_DataOut_6; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_data_7 = DataCorssBarForRead_io_DataOut_7; // @[ShareMem.scala 163:30]
  assign coreRsp_Q_io_enq_bits_activeMask_0 = coreReqActvMask_st2_0; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_1 = coreReqActvMask_st2_1; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_2 = coreReqActvMask_st2_2; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_3 = coreReqActvMask_st2_3; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_4 = coreReqActvMask_st2_4; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_5 = coreReqActvMask_st2_5; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_6 = coreReqActvMask_st2_6; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_enq_bits_activeMask_7 = coreReqActvMask_st2_7; // @[ShareMem.scala 165:36]
  assign coreRsp_Q_io_deq_ready = io_coreRsp_ready; // @[ShareMem.scala 160:20]
  assign DataAccessesRRsp_DataAccess_clock = clock;
  assign DataAccessesRRsp_DataAccess_reset = reset;
  assign DataAccessesRRsp_DataAccess_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_1[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_1[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_1[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_1[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_0_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_1_clock = clock;
  assign DataAccessesRRsp_DataAccess_1_reset = reset;
  assign DataAccessesRRsp_DataAccess_1_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_1_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_3[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_3[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_3[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_3[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_1_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_1_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_2_clock = clock;
  assign DataAccessesRRsp_DataAccess_2_reset = reset;
  assign DataAccessesRRsp_DataAccess_2_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_2_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_5[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_5[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_5[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_5[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_2_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_2_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_3_clock = clock;
  assign DataAccessesRRsp_DataAccess_3_reset = reset;
  assign DataAccessesRRsp_DataAccess_3_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_3_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_7[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_7[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_7[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_7[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_3_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_3_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_4_clock = clock;
  assign DataAccessesRRsp_DataAccess_4_reset = reset;
  assign DataAccessesRRsp_DataAccess_4_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_4_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_9[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_9[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_9[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_9[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_4_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_4_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_5_clock = clock;
  assign DataAccessesRRsp_DataAccess_5_reset = reset;
  assign DataAccessesRRsp_DataAccess_5_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_5_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_11[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_11[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_11[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_11[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_5_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_5_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_6_clock = clock;
  assign DataAccessesRRsp_DataAccess_6_reset = reset;
  assign DataAccessesRRsp_DataAccess_6_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_6_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_13[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_13[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_13[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_13[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_6_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_6_wordOffset1H; // @[ShareMem.scala 139:48]
  assign DataAccessesRRsp_DataAccess_7_clock = clock;
  assign DataAccessesRRsp_DataAccess_7_reset = reset;
  assign DataAccessesRRsp_DataAccess_7_io_r_req_valid = _coreReqisValidWrite_st1_T & _coreReqisValidRead_st1_T_1; // @[ShareMem.scala 142:52]
  assign DataAccessesRRsp_DataAccess_7_io_r_req_bits_setIdx = io_coreReq_bits_setIdx; // @[ShareMem.scala 147:42]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_valid = coreReqisValidWrite_st1; // @[ShareMem.scala 131:31]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_setIdx = coreReq_st1_setIdx; // @[ShareMem.scala 137:39]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_0 = _DataAccessesRRsp_WIRE_15[7:0]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_1 = _DataAccessesRRsp_WIRE_15[15:8]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_2 = _DataAccessesRRsp_WIRE_15[23:16]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_data_3 = _DataAccessesRRsp_WIRE_15[31:24]; // @[ShareMem.scala 132:81]
  assign DataAccessesRRsp_DataAccess_7_io_w_req_bits_waymask = arbAddrCrsbarOut_st1_7_wordOffset1H; // @[ShareMem.scala 139:48]
  always @(posedge clock) begin
    coreReqisValidWrite_st1 <= _coreReqisValidWrite_st1_T & io_coreReq_bits_isWrite; // @[ShareMem.scala 103:59]
    coreReqisValidRead_st1 <= _coreReqisValidWrite_st1_T & ~io_coreReq_bits_isWrite; // @[ShareMem.scala 104:59]
    coreReqisValidRead_st2 <= coreReqisValidRead_st1; // @[ShareMem.scala 105:39]
    coreReqisValidWrite_st2 <= coreReqisValidWrite_st1; // @[ShareMem.scala 106:40]
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_instrId <= io_coreReq_bits_instrId; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_setIdx <= io_coreReq_bits_setIdx; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_0_activeMask <= io_coreReq_bits_perLaneAddr_0_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_1_activeMask <= io_coreReq_bits_perLaneAddr_1_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_2_activeMask <= io_coreReq_bits_perLaneAddr_2_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_3_activeMask <= io_coreReq_bits_perLaneAddr_3_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_4_activeMask <= io_coreReq_bits_perLaneAddr_4_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_5_activeMask <= io_coreReq_bits_perLaneAddr_5_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_6_activeMask <= io_coreReq_bits_perLaneAddr_6_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_perLaneAddr_7_activeMask <= io_coreReq_bits_perLaneAddr_7_activeMask; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_0 <= io_coreReq_bits_data_0; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_1 <= io_coreReq_bits_data_1; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_2 <= io_coreReq_bits_data_2; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_3 <= io_coreReq_bits_data_3; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_4 <= io_coreReq_bits_data_4; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_5 <= io_coreReq_bits_data_5; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_6 <= io_coreReq_bits_data_6; // @[Reg.scala 17:22]
    end
    if (io_coreReq_ready) begin // @[Reg.scala 17:18]
      coreReq_st1_data_7 <= io_coreReq_bits_data_7; // @[Reg.scala 17:22]
    end
    coreReqInstrId_st2 <= coreReq_st1_instrId; // @[ShareMem.scala 109:35]
    coreReqActvMask_st2_0 <= coreReq_st1_perLaneAddr_0_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_1 <= coreReq_st1_perLaneAddr_1_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_2 <= coreReq_st1_perLaneAddr_2_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_3 <= coreReq_st1_perLaneAddr_3_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_4 <= coreReq_st1_perLaneAddr_4_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_5 <= coreReq_st1_perLaneAddr_5_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_6 <= coreReq_st1_perLaneAddr_6_activeMask; // @[ShareMem.scala 110:{44,44}]
    coreReqActvMask_st2_7 <= coreReq_st1_perLaneAddr_7_activeMask; // @[ShareMem.scala 110:{44,44}]
    arbAddrCrsbarOut_st1_0_wordOffset1H <= BankConfArb_io_addrCrsbarOut_0_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_1_wordOffset1H <= BankConfArb_io_addrCrsbarOut_1_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_2_wordOffset1H <= BankConfArb_io_addrCrsbarOut_2_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_3_wordOffset1H <= BankConfArb_io_addrCrsbarOut_3_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_4_wordOffset1H <= BankConfArb_io_addrCrsbarOut_4_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_5_wordOffset1H <= BankConfArb_io_addrCrsbarOut_5_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_6_wordOffset1H <= BankConfArb_io_addrCrsbarOut_6_wordOffset1H; // @[ShareMem.scala 113:37]
    arbAddrCrsbarOut_st1_7_wordOffset1H <= BankConfArb_io_addrCrsbarOut_7_wordOffset1H; // @[ShareMem.scala 113:37]
    arbDataCrsbarSel1H_st1_0 <= BankConfArb_io_dataCrsbarSel1H_0; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_1 <= BankConfArb_io_dataCrsbarSel1H_1; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_2 <= BankConfArb_io_dataCrsbarSel1H_2; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_3 <= BankConfArb_io_dataCrsbarSel1H_3; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_4 <= BankConfArb_io_dataCrsbarSel1H_4; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_5 <= BankConfArb_io_dataCrsbarSel1H_5; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_6 <= BankConfArb_io_dataCrsbarSel1H_6; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st1_7 <= BankConfArb_io_dataCrsbarSel1H_7; // @[ShareMem.scala 114:39]
    arbDataCrsbarSel1H_st2_0 <= arbDataCrsbarSel1H_st1_0; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_1 <= arbDataCrsbarSel1H_st1_1; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_2 <= arbDataCrsbarSel1H_st1_2; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_3 <= arbDataCrsbarSel1H_st1_3; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_4 <= arbDataCrsbarSel1H_st1_4; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_5 <= arbDataCrsbarSel1H_st1_5; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_6 <= arbDataCrsbarSel1H_st1_6; // @[ShareMem.scala 115:39]
    arbDataCrsbarSel1H_st2_7 <= arbDataCrsbarSel1H_st1_7; // @[ShareMem.scala 115:39]
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_0 <= DataAccessesRRsp_0; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_1 <= DataAccessesRRsp_1; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_2 <= DataAccessesRRsp_2; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_3 <= DataAccessesRRsp_3; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_4 <= DataAccessesRRsp_4; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_5 <= DataAccessesRRsp_5; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_6 <= DataAccessesRRsp_6; // @[Reg.scala 17:22]
    end
    if (coreReqisValidRead_st1) begin // @[Reg.scala 17:18]
      dataAccess_data_st2_7 <= DataAccessesRRsp_7; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  coreReqisValidWrite_st1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  coreReqisValidRead_st1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  coreReqisValidRead_st2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  coreReqisValidWrite_st2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  coreReq_st1_instrId = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  coreReq_st1_setIdx = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_0_activeMask = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_1_activeMask = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_2_activeMask = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_3_activeMask = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_4_activeMask = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_5_activeMask = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_6_activeMask = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  coreReq_st1_perLaneAddr_7_activeMask = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  coreReq_st1_data_0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  coreReq_st1_data_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  coreReq_st1_data_2 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  coreReq_st1_data_3 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  coreReq_st1_data_4 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  coreReq_st1_data_5 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  coreReq_st1_data_6 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  coreReq_st1_data_7 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  coreReqInstrId_st2 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  coreReqActvMask_st2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  coreReqActvMask_st2_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  coreReqActvMask_st2_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  coreReqActvMask_st2_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  coreReqActvMask_st2_4 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  coreReqActvMask_st2_5 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  coreReqActvMask_st2_6 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  coreReqActvMask_st2_7 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_0_wordOffset1H = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_1_wordOffset1H = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_2_wordOffset1H = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_3_wordOffset1H = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_4_wordOffset1H = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_5_wordOffset1H = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_6_wordOffset1H = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  arbAddrCrsbarOut_st1_7_wordOffset1H = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_0 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_1 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_2 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_3 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_4 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_5 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_6 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st1_7 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_0 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_1 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_2 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_3 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_4 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_5 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_6 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  arbDataCrsbarSel1H_st2_7 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  dataAccess_data_st2_0 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  dataAccess_data_st2_1 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  dataAccess_data_st2_2 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  dataAccess_data_st2_3 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  dataAccess_data_st2_4 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  dataAccess_data_st2_5 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  dataAccess_data_st2_6 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  dataAccess_data_st2_7 = _RAND_62[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SM_wrapper(
  input         clock,
  input         reset,
  output        io_CTAreq_ready,
  input         io_CTAreq_valid,
  input  [2:0]  io_CTAreq_bits_dispatch2cu_wg_wf_count,
  input  [9:0]  io_CTAreq_bits_dispatch2cu_wf_size_dispatch,
  input  [12:0] io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch,
  input  [12:0] io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch,
  input  [4:0]  io_CTAreq_bits_dispatch2cu_wf_tag_dispatch,
  input  [12:0] io_CTAreq_bits_dispatch2cu_lds_base_dispatch,
  input  [31:0] io_CTAreq_bits_dispatch2cu_start_pc_dispatch,
  output        io_CTArsp_valid,
  output [4:0]  io_CTArsp_bits_cu2dispatch_wf_tag_done,
  output        io_memRsp_ready,
  input         io_memRsp_valid,
  input  [31:0] io_memRsp_bits_d_addr,
  input  [31:0] io_memRsp_bits_d_data_0,
  input  [31:0] io_memRsp_bits_d_data_1,
  input  [31:0] io_memRsp_bits_d_data_2,
  input  [31:0] io_memRsp_bits_d_data_3,
  input  [31:0] io_memRsp_bits_d_data_4,
  input  [31:0] io_memRsp_bits_d_data_5,
  input  [31:0] io_memRsp_bits_d_data_6,
  input  [31:0] io_memRsp_bits_d_data_7,
  input  [2:0]  io_memRsp_bits_d_source,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [2:0]  io_memReq_bits_a_opcode,
  output [31:0] io_memReq_bits_a_addr,
  output [31:0] io_memReq_bits_a_data_0,
  output [31:0] io_memReq_bits_a_data_1,
  output [31:0] io_memReq_bits_a_data_2,
  output [31:0] io_memReq_bits_a_data_3,
  output [31:0] io_memReq_bits_a_data_4,
  output [31:0] io_memReq_bits_a_data_5,
  output [31:0] io_memReq_bits_a_data_6,
  output [31:0] io_memReq_bits_a_data_7,
  output        io_memReq_bits_a_mask_0,
  output        io_memReq_bits_a_mask_1,
  output        io_memReq_bits_a_mask_2,
  output        io_memReq_bits_a_mask_3,
  output        io_memReq_bits_a_mask_4,
  output        io_memReq_bits_a_mask_5,
  output        io_memReq_bits_a_mask_6,
  output        io_memReq_bits_a_mask_7,
  output [2:0]  io_memReq_bits_a_source
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  cta2warp_clock; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_reset; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_io_CTAreq_ready; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_io_CTAreq_valid; // @[GPGPU_top.scala 145:22]
  wire [2:0] cta2warp_io_CTAreq_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 145:22]
  wire [9:0] cta2warp_io_CTAreq_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 145:22]
  wire [12:0] cta2warp_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 145:22]
  wire [12:0] cta2warp_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 145:22]
  wire [4:0] cta2warp_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 145:22]
  wire [12:0] cta2warp_io_CTAreq_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 145:22]
  wire [31:0] cta2warp_io_CTAreq_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_io_CTArsp_valid; // @[GPGPU_top.scala 145:22]
  wire [4:0] cta2warp_io_CTArsp_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_io_warpReq_valid; // @[GPGPU_top.scala 145:22]
  wire [2:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 145:22]
  wire [9:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 145:22]
  wire [12:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 145:22]
  wire [12:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 145:22]
  wire [4:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 145:22]
  wire [12:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 145:22]
  wire [31:0] cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 145:22]
  wire [1:0] cta2warp_io_warpReq_bits_wid; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_io_warpRsp_ready; // @[GPGPU_top.scala 145:22]
  wire  cta2warp_io_warpRsp_valid; // @[GPGPU_top.scala 145:22]
  wire [1:0] cta2warp_io_warpRsp_bits_wid; // @[GPGPU_top.scala 145:22]
  wire [1:0] cta2warp_io_wg_id_lookup; // @[GPGPU_top.scala 145:22]
  wire [4:0] cta2warp_io_wg_id_tag; // @[GPGPU_top.scala 145:22]
  wire  pipe_clock; // @[GPGPU_top.scala 148:18]
  wire  pipe_reset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_icache_req_valid; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_icache_req_bits_addr; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_icache_req_bits_warpid; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_icache_rsp_valid; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_icache_rsp_bits_addr; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_icache_rsp_bits_data; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_icache_rsp_bits_warpid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_icache_rsp_bits_status; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_externalFlushPipe_valid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_externalFlushPipe_bits; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_ready; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_valid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_dcache_req_bits_instrId; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_isWrite; // @[GPGPU_top.scala 148:18]
  wire [21:0] pipe_io_dcache_req_bits_tag; // @[GPGPU_top.scala 148:18]
  wire [4:0] pipe_io_dcache_req_bits_setIdx; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_0_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_0_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_1_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_1_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_2_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_2_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_3_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_3_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_4_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_4_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_5_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_5_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_6_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_6_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_req_bits_perLaneAddr_7_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_dcache_req_bits_perLaneAddr_7_blockOffset; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_0; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_1; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_2; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_3; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_4; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_5; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_6; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_req_bits_data_7; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_ready; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_valid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_dcache_rsp_bits_instrId; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_0; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_1; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_2; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_3; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_4; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_5; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_6; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_dcache_rsp_bits_data_7; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_0; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_1; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_2; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_3; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_4; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_5; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_6; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_dcache_rsp_bits_activeMask_7; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_ready; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_valid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_shared_req_bits_instrId; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_isWrite; // @[GPGPU_top.scala 148:18]
  wire [4:0] pipe_io_shared_req_bits_setIdx; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_0_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_0_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_1_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_1_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_2_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_2_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_3_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_3_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_4_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_4_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_5_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_5_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_6_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_6_blockOffset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_req_bits_perLaneAddr_7_activeMask; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_shared_req_bits_perLaneAddr_7_blockOffset; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_0; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_1; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_2; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_3; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_4; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_5; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_6; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_req_bits_data_7; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_ready; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_valid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_shared_rsp_bits_instrId; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_0; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_1; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_2; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_3; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_4; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_5; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_6; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_shared_rsp_bits_data_7; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_0; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_1; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_2; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_3; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_4; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_5; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_6; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_shared_rsp_bits_activeMask_7; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_pc_reset; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_warpReq_valid; // @[GPGPU_top.scala 148:18]
  wire [2:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 148:18]
  wire [9:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 148:18]
  wire [12:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 148:18]
  wire [12:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 148:18]
  wire [4:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 148:18]
  wire [12:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 148:18]
  wire [31:0] pipe_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_warpReq_bits_wid; // @[GPGPU_top.scala 148:18]
  wire  pipe_io_warpRsp_valid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_warpRsp_bits_wid; // @[GPGPU_top.scala 148:18]
  wire [1:0] pipe_io_wg_id_lookup; // @[GPGPU_top.scala 148:18]
  wire [4:0] pipe_io_wg_id_tag; // @[GPGPU_top.scala 148:18]
  wire  l1Cache2L2Arb_io_memReqVecIn_0_ready; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_0_valid; // @[GPGPU_top.scala 157:29]
  wire [1:0] l1Cache2L2Arb_io_memReqVecIn_0_bits_a_source; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_0_bits_a_addr; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_ready; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_valid; // @[GPGPU_top.scala 157:29]
  wire [2:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_opcode; // @[GPGPU_top.scala 157:29]
  wire [1:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_source; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_addr; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_0; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_1; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_2; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_3; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_4; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_5; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_6; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_7; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_0; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_1; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_2; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_3; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_4; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_5; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_6; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_7; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_ready; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_valid; // @[GPGPU_top.scala 157:29]
  wire [2:0] l1Cache2L2Arb_io_memReqOut_bits_a_opcode; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_addr; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_0; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_1; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_2; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_3; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_4; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_5; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_6; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memReqOut_bits_a_data_7; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_0; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_1; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_2; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_3; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_4; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_5; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_6; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memReqOut_bits_a_mask_7; // @[GPGPU_top.scala 157:29]
  wire [2:0] l1Cache2L2Arb_io_memReqOut_bits_a_source; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memRspIn_ready; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memRspIn_valid; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_addr; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_0; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_1; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_2; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_3; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_4; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_5; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_6; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspIn_bits_d_data_7; // @[GPGPU_top.scala 157:29]
  wire [2:0] l1Cache2L2Arb_io_memRspIn_bits_d_source; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memRspVecOut_0_ready; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memRspVecOut_0_valid; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_addr; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_0; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_1; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_2; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_3; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_4; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_5; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_6; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_7; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memRspVecOut_1_ready; // @[GPGPU_top.scala 157:29]
  wire  l1Cache2L2Arb_io_memRspVecOut_1_valid; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_addr; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_0; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_1; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_2; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_3; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_4; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_5; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_6; // @[GPGPU_top.scala 157:29]
  wire [31:0] l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_7; // @[GPGPU_top.scala 157:29]
  wire  icache_clock; // @[GPGPU_top.scala 161:22]
  wire  icache_reset; // @[GPGPU_top.scala 161:22]
  wire  icache_io_coreReq_ready; // @[GPGPU_top.scala 161:22]
  wire  icache_io_coreReq_valid; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_coreReq_bits_addr; // @[GPGPU_top.scala 161:22]
  wire [1:0] icache_io_coreReq_bits_warpid; // @[GPGPU_top.scala 161:22]
  wire  icache_io_externalFlushPipe_valid; // @[GPGPU_top.scala 161:22]
  wire [1:0] icache_io_externalFlushPipe_bits_warpid; // @[GPGPU_top.scala 161:22]
  wire  icache_io_coreRsp_valid; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_coreRsp_bits_addr; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_coreRsp_bits_data; // @[GPGPU_top.scala 161:22]
  wire [1:0] icache_io_coreRsp_bits_warpid; // @[GPGPU_top.scala 161:22]
  wire [1:0] icache_io_coreRsp_bits_status; // @[GPGPU_top.scala 161:22]
  wire  icache_io_memRsp_ready; // @[GPGPU_top.scala 161:22]
  wire  icache_io_memRsp_valid; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_addr; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_0; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_1; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_2; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_3; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_4; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_5; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_6; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memRsp_bits_d_data_7; // @[GPGPU_top.scala 161:22]
  wire  icache_io_memReq_ready; // @[GPGPU_top.scala 161:22]
  wire  icache_io_memReq_valid; // @[GPGPU_top.scala 161:22]
  wire [1:0] icache_io_memReq_bits_a_source; // @[GPGPU_top.scala 161:22]
  wire [31:0] icache_io_memReq_bits_a_addr; // @[GPGPU_top.scala 161:22]
  wire  dcache_clock; // @[GPGPU_top.scala 196:22]
  wire  dcache_reset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_ready; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_valid; // @[GPGPU_top.scala 196:22]
  wire [1:0] dcache_io_coreReq_bits_instrId; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_isWrite; // @[GPGPU_top.scala 196:22]
  wire [21:0] dcache_io_coreReq_bits_tag; // @[GPGPU_top.scala 196:22]
  wire [4:0] dcache_io_coreReq_bits_setIdx; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_0_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_0_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_1_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_1_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_2_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_2_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_3_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_3_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_4_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_4_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_5_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_5_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_6_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_6_blockOffset; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreReq_bits_perLaneAddr_7_activeMask; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_coreReq_bits_perLaneAddr_7_blockOffset; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_0; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_1; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_2; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_3; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_4; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_5; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_6; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreReq_bits_data_7; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_ready; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_valid; // @[GPGPU_top.scala 196:22]
  wire [1:0] dcache_io_coreRsp_bits_instrId; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_0; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_1; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_2; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_3; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_4; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_5; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_6; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_coreRsp_bits_data_7; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_0; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_1; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_2; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_3; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_4; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_5; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_6; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_coreRsp_bits_activeMask_7; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memRsp_ready; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memRsp_valid; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_addr; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_0; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_1; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_2; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_3; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_4; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_5; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_6; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memRsp_bits_d_data_7; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_ready; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_valid; // @[GPGPU_top.scala 196:22]
  wire [2:0] dcache_io_memReq_bits_a_opcode; // @[GPGPU_top.scala 196:22]
  wire [1:0] dcache_io_memReq_bits_a_source; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_addr; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_0; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_1; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_2; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_3; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_4; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_5; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_6; // @[GPGPU_top.scala 196:22]
  wire [31:0] dcache_io_memReq_bits_a_data_7; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_0; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_1; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_2; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_3; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_4; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_5; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_6; // @[GPGPU_top.scala 196:22]
  wire  dcache_io_memReq_bits_a_mask_7; // @[GPGPU_top.scala 196:22]
  wire  sharedmem_clock; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_reset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_ready; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_valid; // @[GPGPU_top.scala 223:25]
  wire [1:0] sharedmem_io_coreReq_bits_instrId; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_isWrite; // @[GPGPU_top.scala 223:25]
  wire [6:0] sharedmem_io_coreReq_bits_setIdx; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_0_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_0_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_1_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_1_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_2_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_2_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_3_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_3_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_4_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_4_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_5_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_5_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_6_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_6_blockOffset; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreReq_bits_perLaneAddr_7_activeMask; // @[GPGPU_top.scala 223:25]
  wire [2:0] sharedmem_io_coreReq_bits_perLaneAddr_7_blockOffset; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_0; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_1; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_2; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_3; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_4; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_5; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_6; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreReq_bits_data_7; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_ready; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_valid; // @[GPGPU_top.scala 223:25]
  wire [1:0] sharedmem_io_coreRsp_bits_instrId; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_0; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_1; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_2; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_3; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_4; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_5; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_6; // @[GPGPU_top.scala 223:25]
  wire [31:0] sharedmem_io_coreRsp_bits_data_7; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_0; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_1; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_2; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_3; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_4; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_5; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_6; // @[GPGPU_top.scala 223:25]
  wire  sharedmem_io_coreRsp_bits_activeMask_7; // @[GPGPU_top.scala 223:25]
  reg [3:0] value; // @[Counter.scala 62:40]
  wire  wrap = value == 4'h9; // @[Counter.scala 74:24]
  wire [3:0] _value_T_1 = value + 4'h1; // @[Counter.scala 78:24]
  CTA2warp cta2warp ( // @[GPGPU_top.scala 145:22]
    .clock(cta2warp_clock),
    .reset(cta2warp_reset),
    .io_CTAreq_ready(cta2warp_io_CTAreq_ready),
    .io_CTAreq_valid(cta2warp_io_CTAreq_valid),
    .io_CTAreq_bits_dispatch2cu_wg_wf_count(cta2warp_io_CTAreq_bits_dispatch2cu_wg_wf_count),
    .io_CTAreq_bits_dispatch2cu_wf_size_dispatch(cta2warp_io_CTAreq_bits_dispatch2cu_wf_size_dispatch),
    .io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch(cta2warp_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch(cta2warp_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_wf_tag_dispatch(cta2warp_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch),
    .io_CTAreq_bits_dispatch2cu_lds_base_dispatch(cta2warp_io_CTAreq_bits_dispatch2cu_lds_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_start_pc_dispatch(cta2warp_io_CTAreq_bits_dispatch2cu_start_pc_dispatch),
    .io_CTArsp_valid(cta2warp_io_CTArsp_valid),
    .io_CTArsp_bits_cu2dispatch_wf_tag_done(cta2warp_io_CTArsp_bits_cu2dispatch_wf_tag_done),
    .io_warpReq_valid(cta2warp_io_warpReq_valid),
    .io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count(cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch(cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch)
      ,
    .io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(
      cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(
      cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch(cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch(
      cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch(
      cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch),
    .io_warpReq_bits_wid(cta2warp_io_warpReq_bits_wid),
    .io_warpRsp_ready(cta2warp_io_warpRsp_ready),
    .io_warpRsp_valid(cta2warp_io_warpRsp_valid),
    .io_warpRsp_bits_wid(cta2warp_io_warpRsp_bits_wid),
    .io_wg_id_lookup(cta2warp_io_wg_id_lookup),
    .io_wg_id_tag(cta2warp_io_wg_id_tag)
  );
  pipe pipe ( // @[GPGPU_top.scala 148:18]
    .clock(pipe_clock),
    .reset(pipe_reset),
    .io_icache_req_valid(pipe_io_icache_req_valid),
    .io_icache_req_bits_addr(pipe_io_icache_req_bits_addr),
    .io_icache_req_bits_warpid(pipe_io_icache_req_bits_warpid),
    .io_icache_rsp_valid(pipe_io_icache_rsp_valid),
    .io_icache_rsp_bits_addr(pipe_io_icache_rsp_bits_addr),
    .io_icache_rsp_bits_data(pipe_io_icache_rsp_bits_data),
    .io_icache_rsp_bits_warpid(pipe_io_icache_rsp_bits_warpid),
    .io_icache_rsp_bits_status(pipe_io_icache_rsp_bits_status),
    .io_externalFlushPipe_valid(pipe_io_externalFlushPipe_valid),
    .io_externalFlushPipe_bits(pipe_io_externalFlushPipe_bits),
    .io_dcache_req_ready(pipe_io_dcache_req_ready),
    .io_dcache_req_valid(pipe_io_dcache_req_valid),
    .io_dcache_req_bits_instrId(pipe_io_dcache_req_bits_instrId),
    .io_dcache_req_bits_isWrite(pipe_io_dcache_req_bits_isWrite),
    .io_dcache_req_bits_tag(pipe_io_dcache_req_bits_tag),
    .io_dcache_req_bits_setIdx(pipe_io_dcache_req_bits_setIdx),
    .io_dcache_req_bits_perLaneAddr_0_activeMask(pipe_io_dcache_req_bits_perLaneAddr_0_activeMask),
    .io_dcache_req_bits_perLaneAddr_0_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_0_blockOffset),
    .io_dcache_req_bits_perLaneAddr_1_activeMask(pipe_io_dcache_req_bits_perLaneAddr_1_activeMask),
    .io_dcache_req_bits_perLaneAddr_1_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_1_blockOffset),
    .io_dcache_req_bits_perLaneAddr_2_activeMask(pipe_io_dcache_req_bits_perLaneAddr_2_activeMask),
    .io_dcache_req_bits_perLaneAddr_2_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_2_blockOffset),
    .io_dcache_req_bits_perLaneAddr_3_activeMask(pipe_io_dcache_req_bits_perLaneAddr_3_activeMask),
    .io_dcache_req_bits_perLaneAddr_3_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_3_blockOffset),
    .io_dcache_req_bits_perLaneAddr_4_activeMask(pipe_io_dcache_req_bits_perLaneAddr_4_activeMask),
    .io_dcache_req_bits_perLaneAddr_4_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_4_blockOffset),
    .io_dcache_req_bits_perLaneAddr_5_activeMask(pipe_io_dcache_req_bits_perLaneAddr_5_activeMask),
    .io_dcache_req_bits_perLaneAddr_5_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_5_blockOffset),
    .io_dcache_req_bits_perLaneAddr_6_activeMask(pipe_io_dcache_req_bits_perLaneAddr_6_activeMask),
    .io_dcache_req_bits_perLaneAddr_6_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_6_blockOffset),
    .io_dcache_req_bits_perLaneAddr_7_activeMask(pipe_io_dcache_req_bits_perLaneAddr_7_activeMask),
    .io_dcache_req_bits_perLaneAddr_7_blockOffset(pipe_io_dcache_req_bits_perLaneAddr_7_blockOffset),
    .io_dcache_req_bits_data_0(pipe_io_dcache_req_bits_data_0),
    .io_dcache_req_bits_data_1(pipe_io_dcache_req_bits_data_1),
    .io_dcache_req_bits_data_2(pipe_io_dcache_req_bits_data_2),
    .io_dcache_req_bits_data_3(pipe_io_dcache_req_bits_data_3),
    .io_dcache_req_bits_data_4(pipe_io_dcache_req_bits_data_4),
    .io_dcache_req_bits_data_5(pipe_io_dcache_req_bits_data_5),
    .io_dcache_req_bits_data_6(pipe_io_dcache_req_bits_data_6),
    .io_dcache_req_bits_data_7(pipe_io_dcache_req_bits_data_7),
    .io_dcache_rsp_ready(pipe_io_dcache_rsp_ready),
    .io_dcache_rsp_valid(pipe_io_dcache_rsp_valid),
    .io_dcache_rsp_bits_instrId(pipe_io_dcache_rsp_bits_instrId),
    .io_dcache_rsp_bits_data_0(pipe_io_dcache_rsp_bits_data_0),
    .io_dcache_rsp_bits_data_1(pipe_io_dcache_rsp_bits_data_1),
    .io_dcache_rsp_bits_data_2(pipe_io_dcache_rsp_bits_data_2),
    .io_dcache_rsp_bits_data_3(pipe_io_dcache_rsp_bits_data_3),
    .io_dcache_rsp_bits_data_4(pipe_io_dcache_rsp_bits_data_4),
    .io_dcache_rsp_bits_data_5(pipe_io_dcache_rsp_bits_data_5),
    .io_dcache_rsp_bits_data_6(pipe_io_dcache_rsp_bits_data_6),
    .io_dcache_rsp_bits_data_7(pipe_io_dcache_rsp_bits_data_7),
    .io_dcache_rsp_bits_activeMask_0(pipe_io_dcache_rsp_bits_activeMask_0),
    .io_dcache_rsp_bits_activeMask_1(pipe_io_dcache_rsp_bits_activeMask_1),
    .io_dcache_rsp_bits_activeMask_2(pipe_io_dcache_rsp_bits_activeMask_2),
    .io_dcache_rsp_bits_activeMask_3(pipe_io_dcache_rsp_bits_activeMask_3),
    .io_dcache_rsp_bits_activeMask_4(pipe_io_dcache_rsp_bits_activeMask_4),
    .io_dcache_rsp_bits_activeMask_5(pipe_io_dcache_rsp_bits_activeMask_5),
    .io_dcache_rsp_bits_activeMask_6(pipe_io_dcache_rsp_bits_activeMask_6),
    .io_dcache_rsp_bits_activeMask_7(pipe_io_dcache_rsp_bits_activeMask_7),
    .io_shared_req_ready(pipe_io_shared_req_ready),
    .io_shared_req_valid(pipe_io_shared_req_valid),
    .io_shared_req_bits_instrId(pipe_io_shared_req_bits_instrId),
    .io_shared_req_bits_isWrite(pipe_io_shared_req_bits_isWrite),
    .io_shared_req_bits_setIdx(pipe_io_shared_req_bits_setIdx),
    .io_shared_req_bits_perLaneAddr_0_activeMask(pipe_io_shared_req_bits_perLaneAddr_0_activeMask),
    .io_shared_req_bits_perLaneAddr_0_blockOffset(pipe_io_shared_req_bits_perLaneAddr_0_blockOffset),
    .io_shared_req_bits_perLaneAddr_1_activeMask(pipe_io_shared_req_bits_perLaneAddr_1_activeMask),
    .io_shared_req_bits_perLaneAddr_1_blockOffset(pipe_io_shared_req_bits_perLaneAddr_1_blockOffset),
    .io_shared_req_bits_perLaneAddr_2_activeMask(pipe_io_shared_req_bits_perLaneAddr_2_activeMask),
    .io_shared_req_bits_perLaneAddr_2_blockOffset(pipe_io_shared_req_bits_perLaneAddr_2_blockOffset),
    .io_shared_req_bits_perLaneAddr_3_activeMask(pipe_io_shared_req_bits_perLaneAddr_3_activeMask),
    .io_shared_req_bits_perLaneAddr_3_blockOffset(pipe_io_shared_req_bits_perLaneAddr_3_blockOffset),
    .io_shared_req_bits_perLaneAddr_4_activeMask(pipe_io_shared_req_bits_perLaneAddr_4_activeMask),
    .io_shared_req_bits_perLaneAddr_4_blockOffset(pipe_io_shared_req_bits_perLaneAddr_4_blockOffset),
    .io_shared_req_bits_perLaneAddr_5_activeMask(pipe_io_shared_req_bits_perLaneAddr_5_activeMask),
    .io_shared_req_bits_perLaneAddr_5_blockOffset(pipe_io_shared_req_bits_perLaneAddr_5_blockOffset),
    .io_shared_req_bits_perLaneAddr_6_activeMask(pipe_io_shared_req_bits_perLaneAddr_6_activeMask),
    .io_shared_req_bits_perLaneAddr_6_blockOffset(pipe_io_shared_req_bits_perLaneAddr_6_blockOffset),
    .io_shared_req_bits_perLaneAddr_7_activeMask(pipe_io_shared_req_bits_perLaneAddr_7_activeMask),
    .io_shared_req_bits_perLaneAddr_7_blockOffset(pipe_io_shared_req_bits_perLaneAddr_7_blockOffset),
    .io_shared_req_bits_data_0(pipe_io_shared_req_bits_data_0),
    .io_shared_req_bits_data_1(pipe_io_shared_req_bits_data_1),
    .io_shared_req_bits_data_2(pipe_io_shared_req_bits_data_2),
    .io_shared_req_bits_data_3(pipe_io_shared_req_bits_data_3),
    .io_shared_req_bits_data_4(pipe_io_shared_req_bits_data_4),
    .io_shared_req_bits_data_5(pipe_io_shared_req_bits_data_5),
    .io_shared_req_bits_data_6(pipe_io_shared_req_bits_data_6),
    .io_shared_req_bits_data_7(pipe_io_shared_req_bits_data_7),
    .io_shared_rsp_ready(pipe_io_shared_rsp_ready),
    .io_shared_rsp_valid(pipe_io_shared_rsp_valid),
    .io_shared_rsp_bits_instrId(pipe_io_shared_rsp_bits_instrId),
    .io_shared_rsp_bits_data_0(pipe_io_shared_rsp_bits_data_0),
    .io_shared_rsp_bits_data_1(pipe_io_shared_rsp_bits_data_1),
    .io_shared_rsp_bits_data_2(pipe_io_shared_rsp_bits_data_2),
    .io_shared_rsp_bits_data_3(pipe_io_shared_rsp_bits_data_3),
    .io_shared_rsp_bits_data_4(pipe_io_shared_rsp_bits_data_4),
    .io_shared_rsp_bits_data_5(pipe_io_shared_rsp_bits_data_5),
    .io_shared_rsp_bits_data_6(pipe_io_shared_rsp_bits_data_6),
    .io_shared_rsp_bits_data_7(pipe_io_shared_rsp_bits_data_7),
    .io_shared_rsp_bits_activeMask_0(pipe_io_shared_rsp_bits_activeMask_0),
    .io_shared_rsp_bits_activeMask_1(pipe_io_shared_rsp_bits_activeMask_1),
    .io_shared_rsp_bits_activeMask_2(pipe_io_shared_rsp_bits_activeMask_2),
    .io_shared_rsp_bits_activeMask_3(pipe_io_shared_rsp_bits_activeMask_3),
    .io_shared_rsp_bits_activeMask_4(pipe_io_shared_rsp_bits_activeMask_4),
    .io_shared_rsp_bits_activeMask_5(pipe_io_shared_rsp_bits_activeMask_5),
    .io_shared_rsp_bits_activeMask_6(pipe_io_shared_rsp_bits_activeMask_6),
    .io_shared_rsp_bits_activeMask_7(pipe_io_shared_rsp_bits_activeMask_7),
    .io_pc_reset(pipe_io_pc_reset),
    .io_warpReq_valid(pipe_io_warpReq_valid),
    .io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count(pipe_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count),
    .io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch(pipe_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch(pipe_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch)
      ,
    .io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch(pipe_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch)
      ,
    .io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch(pipe_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch(pipe_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch),
    .io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch(pipe_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch),
    .io_warpReq_bits_wid(pipe_io_warpReq_bits_wid),
    .io_warpRsp_valid(pipe_io_warpRsp_valid),
    .io_warpRsp_bits_wid(pipe_io_warpRsp_bits_wid),
    .io_wg_id_lookup(pipe_io_wg_id_lookup),
    .io_wg_id_tag(pipe_io_wg_id_tag)
  );
  L1Cache2L2Arbiter l1Cache2L2Arb ( // @[GPGPU_top.scala 157:29]
    .io_memReqVecIn_0_ready(l1Cache2L2Arb_io_memReqVecIn_0_ready),
    .io_memReqVecIn_0_valid(l1Cache2L2Arb_io_memReqVecIn_0_valid),
    .io_memReqVecIn_0_bits_a_source(l1Cache2L2Arb_io_memReqVecIn_0_bits_a_source),
    .io_memReqVecIn_0_bits_a_addr(l1Cache2L2Arb_io_memReqVecIn_0_bits_a_addr),
    .io_memReqVecIn_1_ready(l1Cache2L2Arb_io_memReqVecIn_1_ready),
    .io_memReqVecIn_1_valid(l1Cache2L2Arb_io_memReqVecIn_1_valid),
    .io_memReqVecIn_1_bits_a_opcode(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_opcode),
    .io_memReqVecIn_1_bits_a_source(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_source),
    .io_memReqVecIn_1_bits_a_addr(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_addr),
    .io_memReqVecIn_1_bits_a_data_0(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_0),
    .io_memReqVecIn_1_bits_a_data_1(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_1),
    .io_memReqVecIn_1_bits_a_data_2(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_2),
    .io_memReqVecIn_1_bits_a_data_3(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_3),
    .io_memReqVecIn_1_bits_a_data_4(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_4),
    .io_memReqVecIn_1_bits_a_data_5(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_5),
    .io_memReqVecIn_1_bits_a_data_6(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_6),
    .io_memReqVecIn_1_bits_a_data_7(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_7),
    .io_memReqVecIn_1_bits_a_mask_0(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_0),
    .io_memReqVecIn_1_bits_a_mask_1(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_1),
    .io_memReqVecIn_1_bits_a_mask_2(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_2),
    .io_memReqVecIn_1_bits_a_mask_3(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_3),
    .io_memReqVecIn_1_bits_a_mask_4(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_4),
    .io_memReqVecIn_1_bits_a_mask_5(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_5),
    .io_memReqVecIn_1_bits_a_mask_6(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_6),
    .io_memReqVecIn_1_bits_a_mask_7(l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_7),
    .io_memReqOut_ready(l1Cache2L2Arb_io_memReqOut_ready),
    .io_memReqOut_valid(l1Cache2L2Arb_io_memReqOut_valid),
    .io_memReqOut_bits_a_opcode(l1Cache2L2Arb_io_memReqOut_bits_a_opcode),
    .io_memReqOut_bits_a_addr(l1Cache2L2Arb_io_memReqOut_bits_a_addr),
    .io_memReqOut_bits_a_data_0(l1Cache2L2Arb_io_memReqOut_bits_a_data_0),
    .io_memReqOut_bits_a_data_1(l1Cache2L2Arb_io_memReqOut_bits_a_data_1),
    .io_memReqOut_bits_a_data_2(l1Cache2L2Arb_io_memReqOut_bits_a_data_2),
    .io_memReqOut_bits_a_data_3(l1Cache2L2Arb_io_memReqOut_bits_a_data_3),
    .io_memReqOut_bits_a_data_4(l1Cache2L2Arb_io_memReqOut_bits_a_data_4),
    .io_memReqOut_bits_a_data_5(l1Cache2L2Arb_io_memReqOut_bits_a_data_5),
    .io_memReqOut_bits_a_data_6(l1Cache2L2Arb_io_memReqOut_bits_a_data_6),
    .io_memReqOut_bits_a_data_7(l1Cache2L2Arb_io_memReqOut_bits_a_data_7),
    .io_memReqOut_bits_a_mask_0(l1Cache2L2Arb_io_memReqOut_bits_a_mask_0),
    .io_memReqOut_bits_a_mask_1(l1Cache2L2Arb_io_memReqOut_bits_a_mask_1),
    .io_memReqOut_bits_a_mask_2(l1Cache2L2Arb_io_memReqOut_bits_a_mask_2),
    .io_memReqOut_bits_a_mask_3(l1Cache2L2Arb_io_memReqOut_bits_a_mask_3),
    .io_memReqOut_bits_a_mask_4(l1Cache2L2Arb_io_memReqOut_bits_a_mask_4),
    .io_memReqOut_bits_a_mask_5(l1Cache2L2Arb_io_memReqOut_bits_a_mask_5),
    .io_memReqOut_bits_a_mask_6(l1Cache2L2Arb_io_memReqOut_bits_a_mask_6),
    .io_memReqOut_bits_a_mask_7(l1Cache2L2Arb_io_memReqOut_bits_a_mask_7),
    .io_memReqOut_bits_a_source(l1Cache2L2Arb_io_memReqOut_bits_a_source),
    .io_memRspIn_ready(l1Cache2L2Arb_io_memRspIn_ready),
    .io_memRspIn_valid(l1Cache2L2Arb_io_memRspIn_valid),
    .io_memRspIn_bits_d_addr(l1Cache2L2Arb_io_memRspIn_bits_d_addr),
    .io_memRspIn_bits_d_data_0(l1Cache2L2Arb_io_memRspIn_bits_d_data_0),
    .io_memRspIn_bits_d_data_1(l1Cache2L2Arb_io_memRspIn_bits_d_data_1),
    .io_memRspIn_bits_d_data_2(l1Cache2L2Arb_io_memRspIn_bits_d_data_2),
    .io_memRspIn_bits_d_data_3(l1Cache2L2Arb_io_memRspIn_bits_d_data_3),
    .io_memRspIn_bits_d_data_4(l1Cache2L2Arb_io_memRspIn_bits_d_data_4),
    .io_memRspIn_bits_d_data_5(l1Cache2L2Arb_io_memRspIn_bits_d_data_5),
    .io_memRspIn_bits_d_data_6(l1Cache2L2Arb_io_memRspIn_bits_d_data_6),
    .io_memRspIn_bits_d_data_7(l1Cache2L2Arb_io_memRspIn_bits_d_data_7),
    .io_memRspIn_bits_d_source(l1Cache2L2Arb_io_memRspIn_bits_d_source),
    .io_memRspVecOut_0_ready(l1Cache2L2Arb_io_memRspVecOut_0_ready),
    .io_memRspVecOut_0_valid(l1Cache2L2Arb_io_memRspVecOut_0_valid),
    .io_memRspVecOut_0_bits_d_addr(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_addr),
    .io_memRspVecOut_0_bits_d_data_0(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_0),
    .io_memRspVecOut_0_bits_d_data_1(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_1),
    .io_memRspVecOut_0_bits_d_data_2(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_2),
    .io_memRspVecOut_0_bits_d_data_3(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_3),
    .io_memRspVecOut_0_bits_d_data_4(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_4),
    .io_memRspVecOut_0_bits_d_data_5(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_5),
    .io_memRspVecOut_0_bits_d_data_6(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_6),
    .io_memRspVecOut_0_bits_d_data_7(l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_7),
    .io_memRspVecOut_1_ready(l1Cache2L2Arb_io_memRspVecOut_1_ready),
    .io_memRspVecOut_1_valid(l1Cache2L2Arb_io_memRspVecOut_1_valid),
    .io_memRspVecOut_1_bits_d_addr(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_addr),
    .io_memRspVecOut_1_bits_d_data_0(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_0),
    .io_memRspVecOut_1_bits_d_data_1(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_1),
    .io_memRspVecOut_1_bits_d_data_2(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_2),
    .io_memRspVecOut_1_bits_d_data_3(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_3),
    .io_memRspVecOut_1_bits_d_data_4(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_4),
    .io_memRspVecOut_1_bits_d_data_5(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_5),
    .io_memRspVecOut_1_bits_d_data_6(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_6),
    .io_memRspVecOut_1_bits_d_data_7(l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_7)
  );
  InstructionCache icache ( // @[GPGPU_top.scala 161:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_coreReq_ready(icache_io_coreReq_ready),
    .io_coreReq_valid(icache_io_coreReq_valid),
    .io_coreReq_bits_addr(icache_io_coreReq_bits_addr),
    .io_coreReq_bits_warpid(icache_io_coreReq_bits_warpid),
    .io_externalFlushPipe_valid(icache_io_externalFlushPipe_valid),
    .io_externalFlushPipe_bits_warpid(icache_io_externalFlushPipe_bits_warpid),
    .io_coreRsp_valid(icache_io_coreRsp_valid),
    .io_coreRsp_bits_addr(icache_io_coreRsp_bits_addr),
    .io_coreRsp_bits_data(icache_io_coreRsp_bits_data),
    .io_coreRsp_bits_warpid(icache_io_coreRsp_bits_warpid),
    .io_coreRsp_bits_status(icache_io_coreRsp_bits_status),
    .io_memRsp_ready(icache_io_memRsp_ready),
    .io_memRsp_valid(icache_io_memRsp_valid),
    .io_memRsp_bits_d_addr(icache_io_memRsp_bits_d_addr),
    .io_memRsp_bits_d_data_0(icache_io_memRsp_bits_d_data_0),
    .io_memRsp_bits_d_data_1(icache_io_memRsp_bits_d_data_1),
    .io_memRsp_bits_d_data_2(icache_io_memRsp_bits_d_data_2),
    .io_memRsp_bits_d_data_3(icache_io_memRsp_bits_d_data_3),
    .io_memRsp_bits_d_data_4(icache_io_memRsp_bits_d_data_4),
    .io_memRsp_bits_d_data_5(icache_io_memRsp_bits_d_data_5),
    .io_memRsp_bits_d_data_6(icache_io_memRsp_bits_d_data_6),
    .io_memRsp_bits_d_data_7(icache_io_memRsp_bits_d_data_7),
    .io_memReq_ready(icache_io_memReq_ready),
    .io_memReq_valid(icache_io_memReq_valid),
    .io_memReq_bits_a_source(icache_io_memReq_bits_a_source),
    .io_memReq_bits_a_addr(icache_io_memReq_bits_a_addr)
  );
  DataCache dcache ( // @[GPGPU_top.scala 196:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_coreReq_ready(dcache_io_coreReq_ready),
    .io_coreReq_valid(dcache_io_coreReq_valid),
    .io_coreReq_bits_instrId(dcache_io_coreReq_bits_instrId),
    .io_coreReq_bits_isWrite(dcache_io_coreReq_bits_isWrite),
    .io_coreReq_bits_tag(dcache_io_coreReq_bits_tag),
    .io_coreReq_bits_setIdx(dcache_io_coreReq_bits_setIdx),
    .io_coreReq_bits_perLaneAddr_0_activeMask(dcache_io_coreReq_bits_perLaneAddr_0_activeMask),
    .io_coreReq_bits_perLaneAddr_0_blockOffset(dcache_io_coreReq_bits_perLaneAddr_0_blockOffset),
    .io_coreReq_bits_perLaneAddr_1_activeMask(dcache_io_coreReq_bits_perLaneAddr_1_activeMask),
    .io_coreReq_bits_perLaneAddr_1_blockOffset(dcache_io_coreReq_bits_perLaneAddr_1_blockOffset),
    .io_coreReq_bits_perLaneAddr_2_activeMask(dcache_io_coreReq_bits_perLaneAddr_2_activeMask),
    .io_coreReq_bits_perLaneAddr_2_blockOffset(dcache_io_coreReq_bits_perLaneAddr_2_blockOffset),
    .io_coreReq_bits_perLaneAddr_3_activeMask(dcache_io_coreReq_bits_perLaneAddr_3_activeMask),
    .io_coreReq_bits_perLaneAddr_3_blockOffset(dcache_io_coreReq_bits_perLaneAddr_3_blockOffset),
    .io_coreReq_bits_perLaneAddr_4_activeMask(dcache_io_coreReq_bits_perLaneAddr_4_activeMask),
    .io_coreReq_bits_perLaneAddr_4_blockOffset(dcache_io_coreReq_bits_perLaneAddr_4_blockOffset),
    .io_coreReq_bits_perLaneAddr_5_activeMask(dcache_io_coreReq_bits_perLaneAddr_5_activeMask),
    .io_coreReq_bits_perLaneAddr_5_blockOffset(dcache_io_coreReq_bits_perLaneAddr_5_blockOffset),
    .io_coreReq_bits_perLaneAddr_6_activeMask(dcache_io_coreReq_bits_perLaneAddr_6_activeMask),
    .io_coreReq_bits_perLaneAddr_6_blockOffset(dcache_io_coreReq_bits_perLaneAddr_6_blockOffset),
    .io_coreReq_bits_perLaneAddr_7_activeMask(dcache_io_coreReq_bits_perLaneAddr_7_activeMask),
    .io_coreReq_bits_perLaneAddr_7_blockOffset(dcache_io_coreReq_bits_perLaneAddr_7_blockOffset),
    .io_coreReq_bits_data_0(dcache_io_coreReq_bits_data_0),
    .io_coreReq_bits_data_1(dcache_io_coreReq_bits_data_1),
    .io_coreReq_bits_data_2(dcache_io_coreReq_bits_data_2),
    .io_coreReq_bits_data_3(dcache_io_coreReq_bits_data_3),
    .io_coreReq_bits_data_4(dcache_io_coreReq_bits_data_4),
    .io_coreReq_bits_data_5(dcache_io_coreReq_bits_data_5),
    .io_coreReq_bits_data_6(dcache_io_coreReq_bits_data_6),
    .io_coreReq_bits_data_7(dcache_io_coreReq_bits_data_7),
    .io_coreRsp_ready(dcache_io_coreRsp_ready),
    .io_coreRsp_valid(dcache_io_coreRsp_valid),
    .io_coreRsp_bits_instrId(dcache_io_coreRsp_bits_instrId),
    .io_coreRsp_bits_data_0(dcache_io_coreRsp_bits_data_0),
    .io_coreRsp_bits_data_1(dcache_io_coreRsp_bits_data_1),
    .io_coreRsp_bits_data_2(dcache_io_coreRsp_bits_data_2),
    .io_coreRsp_bits_data_3(dcache_io_coreRsp_bits_data_3),
    .io_coreRsp_bits_data_4(dcache_io_coreRsp_bits_data_4),
    .io_coreRsp_bits_data_5(dcache_io_coreRsp_bits_data_5),
    .io_coreRsp_bits_data_6(dcache_io_coreRsp_bits_data_6),
    .io_coreRsp_bits_data_7(dcache_io_coreRsp_bits_data_7),
    .io_coreRsp_bits_activeMask_0(dcache_io_coreRsp_bits_activeMask_0),
    .io_coreRsp_bits_activeMask_1(dcache_io_coreRsp_bits_activeMask_1),
    .io_coreRsp_bits_activeMask_2(dcache_io_coreRsp_bits_activeMask_2),
    .io_coreRsp_bits_activeMask_3(dcache_io_coreRsp_bits_activeMask_3),
    .io_coreRsp_bits_activeMask_4(dcache_io_coreRsp_bits_activeMask_4),
    .io_coreRsp_bits_activeMask_5(dcache_io_coreRsp_bits_activeMask_5),
    .io_coreRsp_bits_activeMask_6(dcache_io_coreRsp_bits_activeMask_6),
    .io_coreRsp_bits_activeMask_7(dcache_io_coreRsp_bits_activeMask_7),
    .io_memRsp_ready(dcache_io_memRsp_ready),
    .io_memRsp_valid(dcache_io_memRsp_valid),
    .io_memRsp_bits_d_addr(dcache_io_memRsp_bits_d_addr),
    .io_memRsp_bits_d_data_0(dcache_io_memRsp_bits_d_data_0),
    .io_memRsp_bits_d_data_1(dcache_io_memRsp_bits_d_data_1),
    .io_memRsp_bits_d_data_2(dcache_io_memRsp_bits_d_data_2),
    .io_memRsp_bits_d_data_3(dcache_io_memRsp_bits_d_data_3),
    .io_memRsp_bits_d_data_4(dcache_io_memRsp_bits_d_data_4),
    .io_memRsp_bits_d_data_5(dcache_io_memRsp_bits_d_data_5),
    .io_memRsp_bits_d_data_6(dcache_io_memRsp_bits_d_data_6),
    .io_memRsp_bits_d_data_7(dcache_io_memRsp_bits_d_data_7),
    .io_memReq_ready(dcache_io_memReq_ready),
    .io_memReq_valid(dcache_io_memReq_valid),
    .io_memReq_bits_a_opcode(dcache_io_memReq_bits_a_opcode),
    .io_memReq_bits_a_source(dcache_io_memReq_bits_a_source),
    .io_memReq_bits_a_addr(dcache_io_memReq_bits_a_addr),
    .io_memReq_bits_a_data_0(dcache_io_memReq_bits_a_data_0),
    .io_memReq_bits_a_data_1(dcache_io_memReq_bits_a_data_1),
    .io_memReq_bits_a_data_2(dcache_io_memReq_bits_a_data_2),
    .io_memReq_bits_a_data_3(dcache_io_memReq_bits_a_data_3),
    .io_memReq_bits_a_data_4(dcache_io_memReq_bits_a_data_4),
    .io_memReq_bits_a_data_5(dcache_io_memReq_bits_a_data_5),
    .io_memReq_bits_a_data_6(dcache_io_memReq_bits_a_data_6),
    .io_memReq_bits_a_data_7(dcache_io_memReq_bits_a_data_7),
    .io_memReq_bits_a_mask_0(dcache_io_memReq_bits_a_mask_0),
    .io_memReq_bits_a_mask_1(dcache_io_memReq_bits_a_mask_1),
    .io_memReq_bits_a_mask_2(dcache_io_memReq_bits_a_mask_2),
    .io_memReq_bits_a_mask_3(dcache_io_memReq_bits_a_mask_3),
    .io_memReq_bits_a_mask_4(dcache_io_memReq_bits_a_mask_4),
    .io_memReq_bits_a_mask_5(dcache_io_memReq_bits_a_mask_5),
    .io_memReq_bits_a_mask_6(dcache_io_memReq_bits_a_mask_6),
    .io_memReq_bits_a_mask_7(dcache_io_memReq_bits_a_mask_7)
  );
  SharedMemory sharedmem ( // @[GPGPU_top.scala 223:25]
    .clock(sharedmem_clock),
    .reset(sharedmem_reset),
    .io_coreReq_ready(sharedmem_io_coreReq_ready),
    .io_coreReq_valid(sharedmem_io_coreReq_valid),
    .io_coreReq_bits_instrId(sharedmem_io_coreReq_bits_instrId),
    .io_coreReq_bits_isWrite(sharedmem_io_coreReq_bits_isWrite),
    .io_coreReq_bits_setIdx(sharedmem_io_coreReq_bits_setIdx),
    .io_coreReq_bits_perLaneAddr_0_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_0_activeMask),
    .io_coreReq_bits_perLaneAddr_0_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_0_blockOffset),
    .io_coreReq_bits_perLaneAddr_1_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_1_activeMask),
    .io_coreReq_bits_perLaneAddr_1_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_1_blockOffset),
    .io_coreReq_bits_perLaneAddr_2_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_2_activeMask),
    .io_coreReq_bits_perLaneAddr_2_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_2_blockOffset),
    .io_coreReq_bits_perLaneAddr_3_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_3_activeMask),
    .io_coreReq_bits_perLaneAddr_3_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_3_blockOffset),
    .io_coreReq_bits_perLaneAddr_4_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_4_activeMask),
    .io_coreReq_bits_perLaneAddr_4_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_4_blockOffset),
    .io_coreReq_bits_perLaneAddr_5_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_5_activeMask),
    .io_coreReq_bits_perLaneAddr_5_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_5_blockOffset),
    .io_coreReq_bits_perLaneAddr_6_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_6_activeMask),
    .io_coreReq_bits_perLaneAddr_6_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_6_blockOffset),
    .io_coreReq_bits_perLaneAddr_7_activeMask(sharedmem_io_coreReq_bits_perLaneAddr_7_activeMask),
    .io_coreReq_bits_perLaneAddr_7_blockOffset(sharedmem_io_coreReq_bits_perLaneAddr_7_blockOffset),
    .io_coreReq_bits_data_0(sharedmem_io_coreReq_bits_data_0),
    .io_coreReq_bits_data_1(sharedmem_io_coreReq_bits_data_1),
    .io_coreReq_bits_data_2(sharedmem_io_coreReq_bits_data_2),
    .io_coreReq_bits_data_3(sharedmem_io_coreReq_bits_data_3),
    .io_coreReq_bits_data_4(sharedmem_io_coreReq_bits_data_4),
    .io_coreReq_bits_data_5(sharedmem_io_coreReq_bits_data_5),
    .io_coreReq_bits_data_6(sharedmem_io_coreReq_bits_data_6),
    .io_coreReq_bits_data_7(sharedmem_io_coreReq_bits_data_7),
    .io_coreRsp_ready(sharedmem_io_coreRsp_ready),
    .io_coreRsp_valid(sharedmem_io_coreRsp_valid),
    .io_coreRsp_bits_instrId(sharedmem_io_coreRsp_bits_instrId),
    .io_coreRsp_bits_data_0(sharedmem_io_coreRsp_bits_data_0),
    .io_coreRsp_bits_data_1(sharedmem_io_coreRsp_bits_data_1),
    .io_coreRsp_bits_data_2(sharedmem_io_coreRsp_bits_data_2),
    .io_coreRsp_bits_data_3(sharedmem_io_coreRsp_bits_data_3),
    .io_coreRsp_bits_data_4(sharedmem_io_coreRsp_bits_data_4),
    .io_coreRsp_bits_data_5(sharedmem_io_coreRsp_bits_data_5),
    .io_coreRsp_bits_data_6(sharedmem_io_coreRsp_bits_data_6),
    .io_coreRsp_bits_data_7(sharedmem_io_coreRsp_bits_data_7),
    .io_coreRsp_bits_activeMask_0(sharedmem_io_coreRsp_bits_activeMask_0),
    .io_coreRsp_bits_activeMask_1(sharedmem_io_coreRsp_bits_activeMask_1),
    .io_coreRsp_bits_activeMask_2(sharedmem_io_coreRsp_bits_activeMask_2),
    .io_coreRsp_bits_activeMask_3(sharedmem_io_coreRsp_bits_activeMask_3),
    .io_coreRsp_bits_activeMask_4(sharedmem_io_coreRsp_bits_activeMask_4),
    .io_coreRsp_bits_activeMask_5(sharedmem_io_coreRsp_bits_activeMask_5),
    .io_coreRsp_bits_activeMask_6(sharedmem_io_coreRsp_bits_activeMask_6),
    .io_coreRsp_bits_activeMask_7(sharedmem_io_coreRsp_bits_activeMask_7)
  );
  assign io_CTAreq_ready = cta2warp_io_CTAreq_ready; // @[GPGPU_top.scala 146:21]
  assign io_CTArsp_valid = cta2warp_io_CTArsp_valid; // @[GPGPU_top.scala 147:21]
  assign io_CTArsp_bits_cu2dispatch_wf_tag_done = cta2warp_io_CTArsp_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 147:21]
  assign io_memRsp_ready = l1Cache2L2Arb_io_memRspIn_ready; // @[GPGPU_top.scala 159:29]
  assign io_memReq_valid = l1Cache2L2Arb_io_memReqOut_valid; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_opcode = l1Cache2L2Arb_io_memReqOut_bits_a_opcode; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_addr = l1Cache2L2Arb_io_memReqOut_bits_a_addr; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_0 = l1Cache2L2Arb_io_memReqOut_bits_a_data_0; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_1 = l1Cache2L2Arb_io_memReqOut_bits_a_data_1; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_2 = l1Cache2L2Arb_io_memReqOut_bits_a_data_2; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_3 = l1Cache2L2Arb_io_memReqOut_bits_a_data_3; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_4 = l1Cache2L2Arb_io_memReqOut_bits_a_data_4; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_5 = l1Cache2L2Arb_io_memReqOut_bits_a_data_5; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_6 = l1Cache2L2Arb_io_memReqOut_bits_a_data_6; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_data_7 = l1Cache2L2Arb_io_memReqOut_bits_a_data_7; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_0 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_0; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_1 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_1; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_2 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_2; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_3 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_3; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_4 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_4; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_5 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_5; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_6 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_6; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_mask_7 = l1Cache2L2Arb_io_memReqOut_bits_a_mask_7; // @[GPGPU_top.scala 158:13]
  assign io_memReq_bits_a_source = l1Cache2L2Arb_io_memReqOut_bits_a_source; // @[GPGPU_top.scala 158:13]
  assign cta2warp_clock = clock;
  assign cta2warp_reset = reset;
  assign cta2warp_io_CTAreq_valid = io_CTAreq_valid; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_wg_wf_count = io_CTAreq_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_wf_size_dispatch = io_CTAreq_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch = io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch = io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch = io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_lds_base_dispatch = io_CTAreq_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_CTAreq_bits_dispatch2cu_start_pc_dispatch = io_CTAreq_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 146:21]
  assign cta2warp_io_warpRsp_valid = pipe_io_warpRsp_valid; // @[GPGPU_top.scala 154:18]
  assign cta2warp_io_warpRsp_bits_wid = pipe_io_warpRsp_bits_wid; // @[GPGPU_top.scala 154:18]
  assign cta2warp_io_wg_id_lookup = pipe_io_wg_id_lookup; // @[GPGPU_top.scala 156:27]
  assign pipe_clock = clock;
  assign pipe_reset = reset;
  assign pipe_io_icache_rsp_valid = icache_io_coreRsp_valid; // @[GPGPU_top.scala 186:27]
  assign pipe_io_icache_rsp_bits_addr = icache_io_coreRsp_bits_addr; // @[GPGPU_top.scala 189:31]
  assign pipe_io_icache_rsp_bits_data = icache_io_coreRsp_bits_data; // @[GPGPU_top.scala 188:31]
  assign pipe_io_icache_rsp_bits_warpid = icache_io_coreRsp_bits_warpid; // @[GPGPU_top.scala 187:33]
  assign pipe_io_icache_rsp_bits_status = icache_io_coreRsp_bits_status; // @[GPGPU_top.scala 190:33]
  assign pipe_io_dcache_req_ready = dcache_io_coreReq_ready; // @[GPGPU_top.scala 207:27]
  assign pipe_io_dcache_rsp_valid = dcache_io_coreRsp_valid; // @[GPGPU_top.scala 216:27]
  assign pipe_io_dcache_rsp_bits_instrId = dcache_io_coreRsp_bits_instrId; // @[GPGPU_top.scala 217:34]
  assign pipe_io_dcache_rsp_bits_data_0 = dcache_io_coreRsp_bits_data_0; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_1 = dcache_io_coreRsp_bits_data_1; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_2 = dcache_io_coreRsp_bits_data_2; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_3 = dcache_io_coreRsp_bits_data_3; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_4 = dcache_io_coreRsp_bits_data_4; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_5 = dcache_io_coreRsp_bits_data_5; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_6 = dcache_io_coreRsp_bits_data_6; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_data_7 = dcache_io_coreRsp_bits_data_7; // @[GPGPU_top.scala 218:31]
  assign pipe_io_dcache_rsp_bits_activeMask_0 = dcache_io_coreRsp_bits_activeMask_0; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_1 = dcache_io_coreRsp_bits_activeMask_1; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_2 = dcache_io_coreRsp_bits_activeMask_2; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_3 = dcache_io_coreRsp_bits_activeMask_3; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_4 = dcache_io_coreRsp_bits_activeMask_4; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_5 = dcache_io_coreRsp_bits_activeMask_5; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_6 = dcache_io_coreRsp_bits_activeMask_6; // @[GPGPU_top.scala 219:37]
  assign pipe_io_dcache_rsp_bits_activeMask_7 = dcache_io_coreRsp_bits_activeMask_7; // @[GPGPU_top.scala 219:37]
  assign pipe_io_shared_req_ready = sharedmem_io_coreReq_ready; // @[GPGPU_top.scala 230:27]
  assign pipe_io_shared_rsp_valid = sharedmem_io_coreRsp_valid; // @[GPGPU_top.scala 233:27]
  assign pipe_io_shared_rsp_bits_instrId = sharedmem_io_coreRsp_bits_instrId; // @[GPGPU_top.scala 235:34]
  assign pipe_io_shared_rsp_bits_data_0 = sharedmem_io_coreRsp_bits_data_0; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_1 = sharedmem_io_coreRsp_bits_data_1; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_2 = sharedmem_io_coreRsp_bits_data_2; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_3 = sharedmem_io_coreRsp_bits_data_3; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_4 = sharedmem_io_coreRsp_bits_data_4; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_5 = sharedmem_io_coreRsp_bits_data_5; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_6 = sharedmem_io_coreRsp_bits_data_6; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_data_7 = sharedmem_io_coreRsp_bits_data_7; // @[GPGPU_top.scala 234:31]
  assign pipe_io_shared_rsp_bits_activeMask_0 = sharedmem_io_coreRsp_bits_activeMask_0; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_1 = sharedmem_io_coreRsp_bits_activeMask_1; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_2 = sharedmem_io_coreRsp_bits_activeMask_2; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_3 = sharedmem_io_coreRsp_bits_activeMask_3; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_4 = sharedmem_io_coreRsp_bits_activeMask_4; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_5 = sharedmem_io_coreRsp_bits_activeMask_5; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_6 = sharedmem_io_coreRsp_bits_activeMask_6; // @[GPGPU_top.scala 236:37]
  assign pipe_io_shared_rsp_bits_activeMask_7 = sharedmem_io_coreRsp_bits_activeMask_7; // @[GPGPU_top.scala 236:37]
  assign pipe_io_pc_reset = value == 4'h5 ? 1'h0 : 1'h1; // @[GPGPU_top.scala 149:19 152:{24,41}]
  assign pipe_io_warpReq_valid = cta2warp_io_warpReq_valid; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count = cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wg_wf_count
    ; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch =
    cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch =
    cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch =
    cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch =
    cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch =
    cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch =
    cta2warp_io_warpReq_bits_CTAdata_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 153:18]
  assign pipe_io_warpReq_bits_wid = cta2warp_io_warpReq_bits_wid; // @[GPGPU_top.scala 153:18]
  assign pipe_io_wg_id_tag = cta2warp_io_wg_id_tag; // @[GPGPU_top.scala 155:20]
  assign l1Cache2L2Arb_io_memReqVecIn_0_valid = icache_io_memReq_valid; // @[GPGPU_top.scala 170:41]
  assign l1Cache2L2Arb_io_memReqVecIn_0_bits_a_source = icache_io_memReq_bits_a_source; // @[GPGPU_top.scala 174:49]
  assign l1Cache2L2Arb_io_memReqVecIn_0_bits_a_addr = icache_io_memReq_bits_a_addr; // @[GPGPU_top.scala 173:47]
  assign l1Cache2L2Arb_io_memReqVecIn_1_valid = dcache_io_memReq_valid; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_opcode = dcache_io_memReq_bits_a_opcode; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_source = dcache_io_memReq_bits_a_source; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_addr = dcache_io_memReq_bits_a_addr; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_0 = dcache_io_memReq_bits_a_data_0; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_1 = dcache_io_memReq_bits_a_data_1; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_2 = dcache_io_memReq_bits_a_data_2; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_3 = dcache_io_memReq_bits_a_data_3; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_4 = dcache_io_memReq_bits_a_data_4; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_5 = dcache_io_memReq_bits_a_data_5; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_6 = dcache_io_memReq_bits_a_data_6; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_data_7 = dcache_io_memReq_bits_a_data_7; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_0 = dcache_io_memReq_bits_a_mask_0; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_1 = dcache_io_memReq_bits_a_mask_1; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_2 = dcache_io_memReq_bits_a_mask_2; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_3 = dcache_io_memReq_bits_a_mask_3; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_4 = dcache_io_memReq_bits_a_mask_4; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_5 = dcache_io_memReq_bits_a_mask_5; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_6 = dcache_io_memReq_bits_a_mask_6; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqVecIn_1_bits_a_mask_7 = dcache_io_memReq_bits_a_mask_7; // @[GPGPU_top.scala 205:35]
  assign l1Cache2L2Arb_io_memReqOut_ready = io_memReq_ready; // @[GPGPU_top.scala 158:13]
  assign l1Cache2L2Arb_io_memRspIn_valid = io_memRsp_valid; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_addr = io_memRsp_bits_d_addr; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_0 = io_memRsp_bits_d_data_0; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_1 = io_memRsp_bits_d_data_1; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_2 = io_memRsp_bits_d_data_2; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_3 = io_memRsp_bits_d_data_3; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_4 = io_memRsp_bits_d_data_4; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_5 = io_memRsp_bits_d_data_5; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_6 = io_memRsp_bits_d_data_6; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_data_7 = io_memRsp_bits_d_data_7; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspIn_bits_d_source = io_memRsp_bits_d_source; // @[GPGPU_top.scala 159:29]
  assign l1Cache2L2Arb_io_memRspVecOut_0_ready = icache_io_memRsp_ready; // @[GPGPU_top.scala 167:42]
  assign l1Cache2L2Arb_io_memRspVecOut_1_ready = dcache_io_memRsp_ready; // @[GPGPU_top.scala 202:42]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_coreReq_valid = pipe_io_icache_req_valid; // @[GPGPU_top.scala 181:26]
  assign icache_io_coreReq_bits_addr = pipe_io_icache_req_bits_addr; // @[GPGPU_top.scala 182:30]
  assign icache_io_coreReq_bits_warpid = pipe_io_icache_req_bits_warpid; // @[GPGPU_top.scala 183:32]
  assign icache_io_externalFlushPipe_valid = pipe_io_externalFlushPipe_valid; // @[GPGPU_top.scala 194:37]
  assign icache_io_externalFlushPipe_bits_warpid = pipe_io_externalFlushPipe_bits; // @[GPGPU_top.scala 193:43]
  assign icache_io_memRsp_valid = l1Cache2L2Arb_io_memRspVecOut_0_valid; // @[GPGPU_top.scala 163:26]
  assign icache_io_memRsp_bits_d_addr = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_addr; // @[GPGPU_top.scala 164:32]
  assign icache_io_memRsp_bits_d_data_0 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_0; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_1 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_1; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_2 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_2; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_3 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_3; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_4 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_4; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_5 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_5; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_6 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_6; // @[GPGPU_top.scala 165:32]
  assign icache_io_memRsp_bits_d_data_7 = l1Cache2L2Arb_io_memRspVecOut_0_bits_d_data_7; // @[GPGPU_top.scala 165:32]
  assign icache_io_memReq_ready = l1Cache2L2Arb_io_memReqVecIn_0_ready; // @[GPGPU_top.scala 177:26]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_coreReq_valid = pipe_io_dcache_req_valid; // @[GPGPU_top.scala 208:26]
  assign dcache_io_coreReq_bits_instrId = pipe_io_dcache_req_bits_instrId; // @[GPGPU_top.scala 210:33]
  assign dcache_io_coreReq_bits_isWrite = pipe_io_dcache_req_bits_isWrite; // @[GPGPU_top.scala 212:33]
  assign dcache_io_coreReq_bits_tag = pipe_io_dcache_req_bits_tag; // @[GPGPU_top.scala 214:29]
  assign dcache_io_coreReq_bits_setIdx = pipe_io_dcache_req_bits_setIdx; // @[GPGPU_top.scala 211:32]
  assign dcache_io_coreReq_bits_perLaneAddr_0_activeMask = pipe_io_dcache_req_bits_perLaneAddr_0_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_0_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_0_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_1_activeMask = pipe_io_dcache_req_bits_perLaneAddr_1_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_1_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_1_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_2_activeMask = pipe_io_dcache_req_bits_perLaneAddr_2_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_2_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_2_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_3_activeMask = pipe_io_dcache_req_bits_perLaneAddr_3_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_3_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_3_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_4_activeMask = pipe_io_dcache_req_bits_perLaneAddr_4_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_4_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_4_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_5_activeMask = pipe_io_dcache_req_bits_perLaneAddr_5_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_5_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_5_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_6_activeMask = pipe_io_dcache_req_bits_perLaneAddr_6_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_6_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_6_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_7_activeMask = pipe_io_dcache_req_bits_perLaneAddr_7_activeMask; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_perLaneAddr_7_blockOffset = pipe_io_dcache_req_bits_perLaneAddr_7_blockOffset; // @[GPGPU_top.scala 213:37]
  assign dcache_io_coreReq_bits_data_0 = pipe_io_dcache_req_bits_data_0; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_1 = pipe_io_dcache_req_bits_data_1; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_2 = pipe_io_dcache_req_bits_data_2; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_3 = pipe_io_dcache_req_bits_data_3; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_4 = pipe_io_dcache_req_bits_data_4; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_5 = pipe_io_dcache_req_bits_data_5; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_6 = pipe_io_dcache_req_bits_data_6; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreReq_bits_data_7 = pipe_io_dcache_req_bits_data_7; // @[GPGPU_top.scala 209:30]
  assign dcache_io_coreRsp_ready = pipe_io_dcache_rsp_ready; // @[GPGPU_top.scala 221:26]
  assign dcache_io_memRsp_valid = l1Cache2L2Arb_io_memRspVecOut_1_valid; // @[GPGPU_top.scala 198:26]
  assign dcache_io_memRsp_bits_d_addr = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_addr; // @[GPGPU_top.scala 200:32]
  assign dcache_io_memRsp_bits_d_data_0 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_0; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_1 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_1; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_2 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_2; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_3 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_3; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_4 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_4; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_5 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_5; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_6 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_6; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memRsp_bits_d_data_7 = l1Cache2L2Arb_io_memRspVecOut_1_bits_d_data_7; // @[GPGPU_top.scala 201:32]
  assign dcache_io_memReq_ready = l1Cache2L2Arb_io_memReqVecIn_1_ready; // @[GPGPU_top.scala 205:35]
  assign sharedmem_clock = clock;
  assign sharedmem_reset = reset;
  assign sharedmem_io_coreReq_valid = pipe_io_shared_req_valid; // @[GPGPU_top.scala 229:29]
  assign sharedmem_io_coreReq_bits_instrId = pipe_io_shared_req_bits_instrId; // @[GPGPU_top.scala 225:36]
  assign sharedmem_io_coreReq_bits_isWrite = pipe_io_shared_req_bits_isWrite; // @[GPGPU_top.scala 226:36]
  assign sharedmem_io_coreReq_bits_setIdx = {{2'd0}, pipe_io_shared_req_bits_setIdx}; // @[GPGPU_top.scala 227:35]
  assign sharedmem_io_coreReq_bits_perLaneAddr_0_activeMask = pipe_io_shared_req_bits_perLaneAddr_0_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_0_blockOffset = pipe_io_shared_req_bits_perLaneAddr_0_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_1_activeMask = pipe_io_shared_req_bits_perLaneAddr_1_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_1_blockOffset = pipe_io_shared_req_bits_perLaneAddr_1_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_2_activeMask = pipe_io_shared_req_bits_perLaneAddr_2_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_2_blockOffset = pipe_io_shared_req_bits_perLaneAddr_2_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_3_activeMask = pipe_io_shared_req_bits_perLaneAddr_3_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_3_blockOffset = pipe_io_shared_req_bits_perLaneAddr_3_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_4_activeMask = pipe_io_shared_req_bits_perLaneAddr_4_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_4_blockOffset = pipe_io_shared_req_bits_perLaneAddr_4_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_5_activeMask = pipe_io_shared_req_bits_perLaneAddr_5_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_5_blockOffset = pipe_io_shared_req_bits_perLaneAddr_5_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_6_activeMask = pipe_io_shared_req_bits_perLaneAddr_6_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_6_blockOffset = pipe_io_shared_req_bits_perLaneAddr_6_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_7_activeMask = pipe_io_shared_req_bits_perLaneAddr_7_activeMask; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_perLaneAddr_7_blockOffset = pipe_io_shared_req_bits_perLaneAddr_7_blockOffset; // @[GPGPU_top.scala 228:40]
  assign sharedmem_io_coreReq_bits_data_0 = pipe_io_shared_req_bits_data_0; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_1 = pipe_io_shared_req_bits_data_1; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_2 = pipe_io_shared_req_bits_data_2; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_3 = pipe_io_shared_req_bits_data_3; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_4 = pipe_io_shared_req_bits_data_4; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_5 = pipe_io_shared_req_bits_data_5; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_6 = pipe_io_shared_req_bits_data_6; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreReq_bits_data_7 = pipe_io_shared_req_bits_data_7; // @[GPGPU_top.scala 224:33]
  assign sharedmem_io_coreRsp_ready = pipe_io_shared_rsp_ready; // @[GPGPU_top.scala 232:29]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value <= 4'h0; // @[Counter.scala 62:40]
    end else if (value < 4'h5) begin // @[GPGPU_top.scala 151:22]
      if (wrap) begin // @[Counter.scala 88:20]
        value <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SourceA(
  output         io_req_ready,
  input          io_req_valid,
  input  [2:0]   io_req_bits_opcode,
  input  [3:0]   io_req_bits_source,
  input  [25:0]  io_req_bits_tag,
  input  [4:0]   io_req_bits_offset,
  input  [255:0] io_req_bits_data,
  input  [7:0]   io_req_bits_mask,
  input          io_req_bits_set,
  input          io_a_ready,
  output         io_a_valid,
  output [2:0]   io_a_bits_opcode,
  output [3:0]   io_a_bits_source,
  output [31:0]  io_a_bits_address,
  output [31:0]  io_a_bits_mask,
  output [255:0] io_a_bits_data
);
  wire [26:0] io_a_bits_address_base_hi = {io_req_bits_tag,io_req_bits_set}; // @[Cat.scala 31:58]
  wire [3:0] _io_a_bits_mask_T_9 = io_req_bits_mask[0] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_11 = io_req_bits_mask[1] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_13 = io_req_bits_mask[2] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_15 = io_req_bits_mask[3] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_17 = io_req_bits_mask[4] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_19 = io_req_bits_mask[5] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_21 = io_req_bits_mask[6] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _io_a_bits_mask_T_23 = io_req_bits_mask[7] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [15:0] io_a_bits_mask_lo = {_io_a_bits_mask_T_15,_io_a_bits_mask_T_13,_io_a_bits_mask_T_11,_io_a_bits_mask_T_9}; // @[Cat.scala 31:58]
  wire [15:0] io_a_bits_mask_hi = {_io_a_bits_mask_T_23,_io_a_bits_mask_T_21,_io_a_bits_mask_T_19,_io_a_bits_mask_T_17}; // @[Cat.scala 31:58]
  assign io_req_ready = io_a_ready; // @[SourceA.scala 50:16]
  assign io_a_valid = io_req_valid; // @[SourceA.scala 51:14]
  assign io_a_bits_opcode = io_req_bits_opcode; // @[SourceA.scala 52:21]
  assign io_a_bits_source = io_req_bits_source; // @[SourceA.scala 55:21]
  assign io_a_bits_address = {io_a_bits_address_base_hi,io_req_bits_offset}; // @[Cat.scala 31:58]
  assign io_a_bits_mask = {io_a_bits_mask_hi,io_a_bits_mask_lo}; // @[Cat.scala 31:58]
  assign io_a_bits_data = io_req_bits_data; // @[SourceA.scala 58:21]
endmodule
module SourceD(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [2:0]   io_req_bits_opcode,
  input  [3:0]   io_req_bits_source,
  input  [25:0]  io_req_bits_tag,
  input  [4:0]   io_req_bits_offset,
  input  [1:0]   io_req_bits_put,
  input  [255:0] io_req_bits_data,
  input  [7:0]   io_req_bits_mask,
  input          io_req_bits_set,
  input          io_req_bits_hit,
  input  [1:0]   io_req_bits_way,
  input          io_req_bits_from_mem,
  input          io_d_ready,
  output         io_d_valid,
  output [3:0]   io_d_bits_source,
  output [255:0] io_d_bits_data,
  output [31:0]  io_d_bits_address,
  output         io_pb_pop_valid,
  output [1:0]   io_pb_pop_bits_index,
  input  [255:0] io_pb_beat_data,
  input  [7:0]   io_pb_beat_mask,
  output         io_bs_radr_valid,
  output [1:0]   io_bs_radr_bits_way,
  output         io_bs_radr_bits_set,
  output [7:0]   io_bs_radr_bits_mask,
  input  [255:0] io_bs_rdat_data,
  output         io_bs_wadr_valid,
  output [1:0]   io_bs_wadr_bits_way,
  output         io_bs_wadr_bits_set,
  output [7:0]   io_bs_wadr_bits_mask,
  output [255:0] io_bs_wdat_data,
  input          io_a_ready,
  output         io_a_valid,
  output [3:0]   io_a_bits_source,
  output [25:0]  io_a_bits_tag,
  output [4:0]   io_a_bits_offset,
  output [255:0] io_a_bits_data,
  output [7:0]   io_a_bits_mask,
  output         io_a_bits_set
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  _io_pb_pop_valid_T = io_req_ready & io_req_valid; // @[Decoupled.scala 50:35]
  reg [255:0] pb_beat_reg_data; // @[SourceD.scala 71:26]
  reg [7:0] pb_beat_reg_mask; // @[SourceD.scala 71:26]
  reg [1:0] stateReg; // @[SourceD.scala 74:24]
  reg [2:0] s1_req_reg_opcode; // @[SourceD.scala 78:27]
  reg [3:0] s1_req_reg_source; // @[SourceD.scala 78:27]
  reg [25:0] s1_req_reg_tag; // @[SourceD.scala 78:27]
  reg [4:0] s1_req_reg_offset; // @[SourceD.scala 78:27]
  reg [255:0] s1_req_reg_data; // @[SourceD.scala 78:27]
  reg [7:0] s1_req_reg_mask; // @[SourceD.scala 78:27]
  reg  s1_req_reg_set; // @[SourceD.scala 78:27]
  reg  s1_req_reg_hit; // @[SourceD.scala 78:27]
  reg [1:0] s1_req_reg_way; // @[SourceD.scala 78:27]
  reg  s1_req_reg_from_mem; // @[SourceD.scala 78:27]
  wire  _GEN_0 = _io_pb_pop_valid_T ? io_req_bits_from_mem : s1_req_reg_from_mem; // @[SourceD.scala 79:22 80:15 78:27]
  wire  _GEN_2 = _io_pb_pop_valid_T ? io_req_bits_hit : s1_req_reg_hit; // @[SourceD.scala 79:22 80:15 78:27]
  wire [255:0] _GEN_5 = _io_pb_pop_valid_T ? io_req_bits_data : s1_req_reg_data; // @[SourceD.scala 79:22 80:15 78:27]
  wire [2:0] _GEN_11 = _io_pb_pop_valid_T ? io_req_bits_opcode : s1_req_reg_opcode; // @[SourceD.scala 79:22 80:15 78:27]
  wire [255:0] _GEN_13 = _io_pb_pop_valid_T ? io_pb_beat_data : pb_beat_reg_data; // @[SourceD.scala 79:22 81:16 71:26]
  reg  busy; // @[SourceD.scala 83:21]
  wire  _s1_need_w_T_2 = _GEN_11 == 3'h0 | _GEN_11 == 3'h1; // @[SourceD.scala 87:47]
  wire  s1_need_w = (_GEN_11 == 3'h0 | _GEN_11 == 3'h1) & ~_GEN_0 & _GEN_2; // @[SourceD.scala 87:102]
  wire  s1_need_r = _GEN_11 == 3'h4; // @[SourceD.scala 89:32]
  reg  read_sent_reg; // @[SourceD.scala 95:28]
  wire  read_sent = _io_pb_pop_valid_T ? 1'h0 : read_sent_reg; // @[SourceD.scala 101:20]
  reg  sourceA_sent_reg; // @[SourceD.scala 111:31]
  wire  _T_5 = _s1_need_w_T_2 & io_a_ready; // @[SourceD.scala 112:72]
  wire  sourceA_sent = _io_pb_pop_valid_T ? 1'h0 : sourceA_sent_reg; // @[SourceD.scala 117:23]
  reg  write_sent_reg; // @[SourceD.scala 120:29]
  wire  write_sent = _io_pb_pop_valid_T ? 1'h0 : write_sent_reg; // @[SourceD.scala 126:21]
  wire [1:0] _GEN_21 = io_a_ready ? 2'h3 : 2'h2; // @[SourceD.scala 140:30]
  wire [1:0] _GEN_23 = _s1_need_w_T_2 ? _GEN_21 : stateReg; // @[SourceD.scala 139:85 74:24]
  wire  _GEN_26 = s1_need_r | _s1_need_w_T_2; // @[SourceD.scala 136:46 138:16]
  wire  _GEN_28 = _io_pb_pop_valid_T & _GEN_26; // @[SourceD.scala 134:11 135:28]
  wire [1:0] _GEN_30 = io_a_ready ? 2'h3 : stateReg; // @[SourceD.scala 165:23 166:17 74:24]
  wire  _GEN_31 = io_d_ready ? 1'h0 : busy; // @[SourceD.scala 170:24 171:14 83:21]
  wire [1:0] _GEN_32 = io_d_ready ? 2'h0 : stateReg; // @[SourceD.scala 170:24 172:18 74:24]
  wire  _GEN_33 = 2'h3 == stateReg ? _GEN_31 : busy; // @[SourceD.scala 132:19 83:21]
  wire [1:0] _GEN_34 = 2'h3 == stateReg ? _GEN_32 : stateReg; // @[SourceD.scala 132:19 74:24]
  reg [2:0] s_final_req_opcode; // @[SourceD.scala 182:26]
  reg [3:0] s_final_req_source; // @[SourceD.scala 182:26]
  reg [25:0] s_final_req_tag; // @[SourceD.scala 182:26]
  reg [4:0] s_final_req_offset; // @[SourceD.scala 182:26]
  reg  s_final_req_set; // @[SourceD.scala 182:26]
  reg  io_d_valid_REG; // @[SourceD.scala 184:30]
  wire  _io_d_bits_opcode_T = s_final_req_opcode == 3'h4; // @[SourceD.scala 186:45]
  wire [26:0] io_d_bits_address_base_hi = {s_final_req_tag,s_final_req_set}; // @[Cat.scala 31:58]
  assign io_req_ready = ~busy; // @[SourceD.scala 108:20]
  assign io_d_valid = io_d_valid_REG; // @[SourceD.scala 184:21]
  assign io_d_bits_source = s_final_req_source; // @[SourceD.scala 185:21]
  assign io_d_bits_data = _io_d_bits_opcode_T ? io_bs_rdat_data : 256'h0; // @[SourceD.scala 188:26]
  assign io_d_bits_address = {io_d_bits_address_base_hi,s_final_req_offset}; // @[Cat.scala 31:58]
  assign io_pb_pop_valid = _io_pb_pop_valid_T & (io_req_bits_opcode == 3'h0 | io_req_bits_opcode == 3'h1) & ~
    io_req_bits_from_mem & io_req_bits_hit; // @[SourceD.scala 68:137]
  assign io_pb_pop_bits_index = io_req_bits_put; // @[SourceD.scala 69:23]
  assign io_bs_radr_valid = s1_need_r & ~read_sent; // @[SourceD.scala 102:37]
  assign io_bs_radr_bits_way = _io_pb_pop_valid_T ? io_req_bits_way : s1_req_reg_way; // @[SourceD.scala 86:18]
  assign io_bs_radr_bits_set = _io_pb_pop_valid_T ? io_req_bits_set : s1_req_reg_set; // @[SourceD.scala 86:18]
  assign io_bs_radr_bits_mask = _io_pb_pop_valid_T ? io_req_bits_mask : s1_req_reg_mask; // @[SourceD.scala 86:18]
  assign io_bs_wadr_valid = s1_need_w & ~write_sent; // @[SourceD.scala 177:39]
  assign io_bs_wadr_bits_way = _io_pb_pop_valid_T ? io_req_bits_way : s1_req_reg_way; // @[SourceD.scala 86:18]
  assign io_bs_wadr_bits_set = _io_pb_pop_valid_T ? io_req_bits_set : s1_req_reg_set; // @[SourceD.scala 86:18]
  assign io_bs_wadr_bits_mask = _io_pb_pop_valid_T ? io_pb_beat_mask : pb_beat_reg_mask; // @[SourceD.scala 85:19]
  assign io_bs_wdat_data = _io_pb_pop_valid_T ? io_pb_beat_data : pb_beat_reg_data; // @[SourceD.scala 85:19]
  assign io_a_valid = _s1_need_w_T_2 & ~sourceA_sent; // @[SourceD.scala 193:86]
  assign io_a_bits_source = _io_pb_pop_valid_T ? io_req_bits_source : s1_req_reg_source; // @[SourceD.scala 86:18]
  assign io_a_bits_tag = _io_pb_pop_valid_T ? io_req_bits_tag : s1_req_reg_tag; // @[SourceD.scala 86:18]
  assign io_a_bits_offset = _io_pb_pop_valid_T ? io_req_bits_offset : s1_req_reg_offset; // @[SourceD.scala 86:18]
  assign io_a_bits_data = _s1_need_w_T_2 ? _GEN_5 : _GEN_13; // @[SourceD.scala 196:25]
  assign io_a_bits_mask = _io_pb_pop_valid_T ? io_req_bits_mask : s1_req_reg_mask; // @[SourceD.scala 86:18]
  assign io_a_bits_set = _io_pb_pop_valid_T ? io_req_bits_set : s1_req_reg_set; // @[SourceD.scala 86:18]
  always @(posedge clock) begin
    if (reset) begin // @[SourceD.scala 71:26]
      pb_beat_reg_data <= 256'h0; // @[SourceD.scala 71:26]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      pb_beat_reg_data <= io_pb_beat_data; // @[SourceD.scala 81:16]
    end
    if (reset) begin // @[SourceD.scala 71:26]
      pb_beat_reg_mask <= 8'h0; // @[SourceD.scala 71:26]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      pb_beat_reg_mask <= io_pb_beat_mask; // @[SourceD.scala 81:16]
    end
    if (reset) begin // @[SourceD.scala 74:24]
      stateReg <= 2'h0; // @[SourceD.scala 74:24]
    end else if (2'h0 == stateReg) begin // @[SourceD.scala 132:19]
      if (_io_pb_pop_valid_T) begin // @[SourceD.scala 135:28]
        if (s1_need_r) begin // @[SourceD.scala 136:46]
          stateReg <= 2'h3; // @[SourceD.scala 137:20]
        end else begin
          stateReg <= _GEN_23;
        end
      end
    end else if (2'h1 == stateReg) begin // @[SourceD.scala 132:19]
      stateReg <= 2'h3;
    end else if (2'h2 == stateReg) begin // @[SourceD.scala 132:19]
      stateReg <= _GEN_30;
    end else begin
      stateReg <= _GEN_34;
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_opcode <= 3'h5; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_opcode <= io_req_bits_opcode; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_source <= 4'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_source <= io_req_bits_source; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_tag <= 26'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_tag <= io_req_bits_tag; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_offset <= 5'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_offset <= io_req_bits_offset; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_data <= 256'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_data <= io_req_bits_data; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_mask <= 8'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_mask <= io_req_bits_mask; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_set <= 1'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_set <= io_req_bits_set; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_hit <= 1'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_hit <= io_req_bits_hit; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_way <= 2'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_way <= io_req_bits_way; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 78:27]
      s1_req_reg_from_mem <= 1'h0; // @[SourceD.scala 78:27]
    end else if (_io_pb_pop_valid_T) begin // @[SourceD.scala 79:22]
      s1_req_reg_from_mem <= io_req_bits_from_mem; // @[SourceD.scala 80:15]
    end
    if (reset) begin // @[SourceD.scala 83:21]
      busy <= 1'h0; // @[SourceD.scala 83:21]
    end else if (2'h0 == stateReg) begin // @[SourceD.scala 132:19]
      busy <= _GEN_28;
    end else if (!(2'h1 == stateReg)) begin // @[SourceD.scala 132:19]
      if (!(2'h2 == stateReg)) begin // @[SourceD.scala 132:19]
        busy <= _GEN_33;
      end
    end
    if (reset) begin // @[SourceD.scala 95:28]
      read_sent_reg <= 1'h0; // @[SourceD.scala 95:28]
    end else begin
      read_sent_reg <= s1_need_r;
    end
    if (reset) begin // @[SourceD.scala 111:31]
      sourceA_sent_reg <= 1'h0; // @[SourceD.scala 111:31]
    end else begin
      sourceA_sent_reg <= _T_5;
    end
    if (reset) begin // @[SourceD.scala 120:29]
      write_sent_reg <= 1'h0; // @[SourceD.scala 120:29]
    end else begin
      write_sent_reg <= s1_need_w;
    end
    if (_io_pb_pop_valid_T) begin // @[SourceD.scala 86:18]
      s_final_req_opcode <= io_req_bits_opcode;
    end else begin
      s_final_req_opcode <= s1_req_reg_opcode;
    end
    if (_io_pb_pop_valid_T) begin // @[SourceD.scala 86:18]
      s_final_req_source <= io_req_bits_source;
    end else begin
      s_final_req_source <= s1_req_reg_source;
    end
    if (_io_pb_pop_valid_T) begin // @[SourceD.scala 86:18]
      s_final_req_tag <= io_req_bits_tag;
    end else begin
      s_final_req_tag <= s1_req_reg_tag;
    end
    if (_io_pb_pop_valid_T) begin // @[SourceD.scala 86:18]
      s_final_req_offset <= io_req_bits_offset;
    end else begin
      s_final_req_offset <= s1_req_reg_offset;
    end
    if (_io_pb_pop_valid_T) begin // @[SourceD.scala 86:18]
      s_final_req_set <= io_req_bits_set;
    end else begin
      s_final_req_set <= s1_req_reg_set;
    end
    io_d_valid_REG <= stateReg == 2'h3 & s1_need_r; // @[SourceD.scala 184:50]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  pb_beat_reg_data = _RAND_0[255:0];
  _RAND_1 = {1{`RANDOM}};
  pb_beat_reg_mask = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  stateReg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  s1_req_reg_opcode = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  s1_req_reg_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  s1_req_reg_tag = _RAND_5[25:0];
  _RAND_6 = {1{`RANDOM}};
  s1_req_reg_offset = _RAND_6[4:0];
  _RAND_7 = {8{`RANDOM}};
  s1_req_reg_data = _RAND_7[255:0];
  _RAND_8 = {1{`RANDOM}};
  s1_req_reg_mask = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  s1_req_reg_set = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  s1_req_reg_hit = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s1_req_reg_way = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  s1_req_reg_from_mem = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  busy = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  read_sent_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sourceA_sent_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  write_sent_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s_final_req_opcode = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  s_final_req_source = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  s_final_req_tag = _RAND_19[25:0];
  _RAND_20 = {1{`RANDOM}};
  s_final_req_offset = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  s_final_req_set = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  io_d_valid_REG = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ListBuffer(
  input          clock,
  input          reset,
  output         io_push_ready,
  input          io_push_valid,
  input  [1:0]   io_push_bits_index,
  input  [255:0] io_push_bits_data_data,
  input  [7:0]   io_push_bits_data_mask,
  output [3:0]   io_valid,
  input          io_pop_valid,
  input  [1:0]   io_pop_bits,
  output [255:0] io_data_data,
  output [7:0]   io_data_mask,
  input          io_pop2_valid,
  input  [1:0]   io_pop2_bits,
  output [255:0] io_data2_data,
  output [7:0]   io_data2_mask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [287:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] head [0:3]; // @[ListBuffer.scala 51:18]
  wire  head_pop_head_en; // @[ListBuffer.scala 51:18]
  wire [1:0] head_pop_head_addr; // @[ListBuffer.scala 51:18]
  wire [1:0] head_pop_head_data; // @[ListBuffer.scala 51:18]
  wire  head_pop_head2_MPORT_en; // @[ListBuffer.scala 51:18]
  wire [1:0] head_pop_head2_MPORT_addr; // @[ListBuffer.scala 51:18]
  wire [1:0] head_pop_head2_MPORT_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_2_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_2_addr; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_2_mask; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_2_en; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_6_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_6_addr; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_6_mask; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_6_en; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_9_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_9_addr; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_9_mask; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_9_en; // @[ListBuffer.scala 51:18]
  reg [1:0] tail [0:3]; // @[ListBuffer.scala 52:18]
  wire  tail_push_tail_en; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_push_tail_addr; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_push_tail_data; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_4_en; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_4_addr; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_4_data; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_7_en; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_7_addr; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_7_data; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_3_data; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_3_addr; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_3_mask; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_3_en; // @[ListBuffer.scala 52:18]
  reg [1:0] next [0:3]; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_5_en; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_5_addr; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_5_data; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_8_en; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_8_addr; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_8_data; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_1_data; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_1_addr; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_1_mask; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_1_en; // @[ListBuffer.scala 54:18]
  reg [263:0] data [0:3]; // @[ListBuffer.scala 55:18]
  wire  data_io_data2_MPORT_en; // @[ListBuffer.scala 55:18]
  wire [1:0] data_io_data2_MPORT_addr; // @[ListBuffer.scala 55:18]
  wire [263:0] data_io_data2_MPORT_data; // @[ListBuffer.scala 55:18]
  wire  data_io_data_MPORT_en; // @[ListBuffer.scala 55:18]
  wire [1:0] data_io_data_MPORT_addr; // @[ListBuffer.scala 55:18]
  wire [263:0] data_io_data_MPORT_data; // @[ListBuffer.scala 55:18]
  wire [263:0] data_MPORT_data; // @[ListBuffer.scala 55:18]
  wire [1:0] data_MPORT_addr; // @[ListBuffer.scala 55:18]
  wire  data_MPORT_mask; // @[ListBuffer.scala 55:18]
  wire  data_MPORT_en; // @[ListBuffer.scala 55:18]
  reg [3:0] valid; // @[ListBuffer.scala 50:22]
  reg [3:0] used; // @[ListBuffer.scala 53:22]
  wire [3:0] _freeOH_T = ~used; // @[ListBuffer.scala 57:27]
  wire [4:0] _freeOH_T_1 = {_freeOH_T, 1'h0}; // @[package.scala 244:48]
  wire [3:0] _freeOH_T_3 = _freeOH_T | _freeOH_T_1[3:0]; // @[package.scala 244:43]
  wire [5:0] _freeOH_T_4 = {_freeOH_T_3, 2'h0}; // @[package.scala 244:48]
  wire [3:0] _freeOH_T_6 = _freeOH_T_3 | _freeOH_T_4[3:0]; // @[package.scala 244:43]
  wire [4:0] _freeOH_T_8 = {_freeOH_T_6, 1'h0}; // @[ListBuffer.scala 57:44]
  wire [4:0] _freeOH_T_9 = ~_freeOH_T_8; // @[ListBuffer.scala 57:17]
  wire [4:0] _GEN_49 = {{1'd0}, _freeOH_T}; // @[ListBuffer.scala 57:60]
  wire [4:0] freeOH = _freeOH_T_9 & _GEN_49; // @[ListBuffer.scala 57:60]
  wire  freeIdx_hi = freeOH[4]; // @[OneHot.scala 30:18]
  wire [3:0] freeIdx_lo = freeOH[3:0]; // @[OneHot.scala 31:18]
  wire  _freeIdx_T = |freeIdx_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_50 = {{3'd0}, freeIdx_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _freeIdx_T_1 = _GEN_50 | freeIdx_lo; // @[OneHot.scala 32:28]
  wire [1:0] freeIdx_hi_1 = _freeIdx_T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] freeIdx_lo_1 = _freeIdx_T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _freeIdx_T_2 = |freeIdx_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _freeIdx_T_3 = freeIdx_hi_1 | freeIdx_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] freeIdx = {_freeIdx_T,_freeIdx_T_2,_freeIdx_T_3[1]}; // @[Cat.scala 31:58]
  wire [3:0] _push_valid_T = valid >> io_push_bits_index; // @[ListBuffer.scala 70:25]
  wire  push_valid = _push_valid_T[0]; // @[ListBuffer.scala 70:25]
  wire  _T = io_push_ready & io_push_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _valid_set_T = 4'h1 << io_push_bits_index; // @[OneHot.scala 64:12]
  wire  _GEN_7 = push_valid ? 1'h0 : 1'h1; // @[ListBuffer.scala 51:18 77:23]
  wire [3:0] valid_set = _T ? _valid_set_T : 4'h0; // @[ListBuffer.scala 73:25 74:15]
  wire [4:0] _GEN_11 = _T ? freeOH : 5'h0; // @[ListBuffer.scala 73:25 75:14]
  wire  _GEN_19 = _T & push_valid; // @[ListBuffer.scala 54:18 73:25]
  wire [263:0] _io_data2_WIRE_1 = data_io_data2_MPORT_data;
  wire [263:0] _io_data_WIRE_1 = data_io_data_MPORT_data;
  wire [3:0] _T_4 = io_valid >> io_pop_bits; // @[ListBuffer.scala 101:39]
  wire  _T_8 = ~reset; // @[ListBuffer.scala 101:10]
  wire [3:0] _T_11 = io_valid >> io_pop2_bits; // @[ListBuffer.scala 103:43]
  wire [1:0] used_clr_shiftAmount = head_pop_head_data; // @[OneHot.scala 63:49]
  wire [3:0] _used_clr_T = 4'h1 << used_clr_shiftAmount; // @[OneHot.scala 64:12]
  wire [3:0] _valid_clr_T = 4'h1 << io_pop_bits; // @[OneHot.scala 64:12]
  wire [3:0] _GEN_29 = head_pop_head_data == tail_MPORT_4_data ? _valid_clr_T : 4'h0; // @[ListBuffer.scala 108:48 109:17]
  wire [2:0] _T_22 = _GEN_19 & tail_push_tail_data == head_pop_head_data ? freeIdx : {{1'd0}, next_MPORT_5_data}; // @[ListBuffer.scala 111:32]
  wire [3:0] used_clr = io_pop_valid ? _used_clr_T : 4'h0; // @[ListBuffer.scala 106:24 107:14]
  wire [3:0] valid_clr = io_pop_valid ? _GEN_29 : 4'h0; // @[ListBuffer.scala 106:24]
  wire [1:0] pop_head2 = head_pop_head2_MPORT_data;
  wire [3:0] _used_clr_2_T = 4'h1 << pop_head2; // @[OneHot.scala 64:12]
  wire [3:0] _valid_clr_2_T = 4'h1 << io_pop2_bits; // @[OneHot.scala 64:12]
  wire [3:0] _GEN_38 = pop_head2 == tail_MPORT_7_data ? _valid_clr_2_T : 4'h0; // @[ListBuffer.scala 116:55 117:21]
  wire [2:0] _T_28 = _GEN_19 & tail_push_tail_data == pop_head2 ? freeIdx : {{1'd0}, next_MPORT_8_data}; // @[ListBuffer.scala 119:39]
  wire [3:0] used_clr_2 = io_pop2_valid ? _used_clr_2_T : 4'h0; // @[ListBuffer.scala 114:30 115:18]
  wire [3:0] valid_clr_2 = io_pop2_valid ? _GEN_38 : 4'h0; // @[ListBuffer.scala 114:30]
  wire [3:0] _used_T = ~used_clr; // @[ListBuffer.scala 124:24]
  wire [3:0] _used_T_1 = used & _used_T; // @[ListBuffer.scala 124:21]
  wire [3:0] _used_T_2 = ~used_clr_2; // @[ListBuffer.scala 124:46]
  wire [3:0] _used_T_3 = _used_T_1 & _used_T_2; // @[ListBuffer.scala 124:44]
  wire [3:0] used_set = _GEN_11[3:0];
  wire [3:0] _used_T_4 = _used_T_3 | used_set; // @[ListBuffer.scala 124:70]
  wire [3:0] _valid_T = ~valid_clr; // @[ListBuffer.scala 125:24]
  wire [3:0] _valid_T_1 = valid & _valid_T; // @[ListBuffer.scala 125:21]
  wire [3:0] _valid_T_2 = ~valid_clr_2; // @[ListBuffer.scala 125:46]
  wire [3:0] _valid_T_3 = _valid_T_1 & _valid_T_2; // @[ListBuffer.scala 125:44]
  wire [3:0] _valid_T_4 = _valid_T_3 | valid_set; // @[ListBuffer.scala 125:71]
  assign head_pop_head_en = 1'h1;
  assign head_pop_head_addr = io_pop_bits;
  assign head_pop_head_data = head[head_pop_head_addr]; // @[ListBuffer.scala 51:18]
  assign head_pop_head2_MPORT_en = 1'h1;
  assign head_pop_head2_MPORT_addr = io_pop2_bits;
  assign head_pop_head2_MPORT_data = head[head_pop_head2_MPORT_addr]; // @[ListBuffer.scala 51:18]
  assign head_MPORT_2_data = freeIdx[1:0];
  assign head_MPORT_2_addr = io_push_bits_index;
  assign head_MPORT_2_mask = 1'h1;
  assign head_MPORT_2_en = _T & _GEN_7;
  assign head_MPORT_6_data = _T_22[1:0];
  assign head_MPORT_6_addr = io_pop_bits;
  assign head_MPORT_6_mask = 1'h1;
  assign head_MPORT_6_en = io_pop_valid;
  assign head_MPORT_9_data = _T_28[1:0];
  assign head_MPORT_9_addr = io_pop2_bits;
  assign head_MPORT_9_mask = 1'h1;
  assign head_MPORT_9_en = io_pop2_valid;
  assign tail_push_tail_en = 1'h1;
  assign tail_push_tail_addr = io_push_bits_index;
  assign tail_push_tail_data = tail[tail_push_tail_addr]; // @[ListBuffer.scala 52:18]
  assign tail_MPORT_4_en = io_pop_valid;
  assign tail_MPORT_4_addr = io_pop_bits;
  assign tail_MPORT_4_data = tail[tail_MPORT_4_addr]; // @[ListBuffer.scala 52:18]
  assign tail_MPORT_7_en = io_pop2_valid;
  assign tail_MPORT_7_addr = io_pop2_bits;
  assign tail_MPORT_7_data = tail[tail_MPORT_7_addr]; // @[ListBuffer.scala 52:18]
  assign tail_MPORT_3_data = freeIdx[1:0];
  assign tail_MPORT_3_addr = io_push_bits_index;
  assign tail_MPORT_3_mask = 1'h1;
  assign tail_MPORT_3_en = io_push_ready & io_push_valid;
  assign next_MPORT_5_en = io_pop_valid;
  assign next_MPORT_5_addr = head_pop_head_data;
  assign next_MPORT_5_data = next[next_MPORT_5_addr]; // @[ListBuffer.scala 54:18]
  assign next_MPORT_8_en = io_pop2_valid;
  assign next_MPORT_8_addr = head_pop_head2_MPORT_data;
  assign next_MPORT_8_data = next[next_MPORT_8_addr]; // @[ListBuffer.scala 54:18]
  assign next_MPORT_1_data = freeIdx[1:0];
  assign next_MPORT_1_addr = tail_push_tail_data;
  assign next_MPORT_1_mask = 1'h1;
  assign next_MPORT_1_en = _T & push_valid;
  assign data_io_data2_MPORT_en = 1'h1;
  assign data_io_data2_MPORT_addr = head_pop_head2_MPORT_data;
  assign data_io_data2_MPORT_data = data[data_io_data2_MPORT_addr]; // @[ListBuffer.scala 55:18]
  assign data_io_data_MPORT_en = 1'h1;
  assign data_io_data_MPORT_addr = head_pop_head_data;
  assign data_io_data_MPORT_data = data[data_io_data_MPORT_addr]; // @[ListBuffer.scala 55:18]
  assign data_MPORT_data = {io_push_bits_data_data,io_push_bits_data_mask};
  assign data_MPORT_addr = freeIdx[1:0];
  assign data_MPORT_mask = 1'h1;
  assign data_MPORT_en = io_push_ready & io_push_valid;
  assign io_push_ready = ~(&used); // @[ListBuffer.scala 72:20]
  assign io_valid = valid; // @[ListBuffer.scala 98:12]
  assign io_data_data = _io_data_WIRE_1[263:8]; // @[ListBuffer.scala 96:63]
  assign io_data_mask = _io_data_WIRE_1[7:0]; // @[ListBuffer.scala 96:63]
  assign io_data2_data = _io_data2_WIRE_1[263:8]; // @[ListBuffer.scala 92:71]
  assign io_data2_mask = _io_data2_WIRE_1[7:0]; // @[ListBuffer.scala 92:71]
  always @(posedge clock) begin
    if (head_MPORT_2_en & head_MPORT_2_mask) begin
      head[head_MPORT_2_addr] <= head_MPORT_2_data; // @[ListBuffer.scala 51:18]
    end
    if (head_MPORT_6_en & head_MPORT_6_mask) begin
      head[head_MPORT_6_addr] <= head_MPORT_6_data; // @[ListBuffer.scala 51:18]
    end
    if (head_MPORT_9_en & head_MPORT_9_mask) begin
      head[head_MPORT_9_addr] <= head_MPORT_9_data; // @[ListBuffer.scala 51:18]
    end
    if (tail_MPORT_3_en & tail_MPORT_3_mask) begin
      tail[tail_MPORT_3_addr] <= tail_MPORT_3_data; // @[ListBuffer.scala 52:18]
    end
    if (next_MPORT_1_en & next_MPORT_1_mask) begin
      next[next_MPORT_1_addr] <= next_MPORT_1_data; // @[ListBuffer.scala 54:18]
    end
    if (data_MPORT_en & data_MPORT_mask) begin
      data[data_MPORT_addr] <= data_MPORT_data; // @[ListBuffer.scala 55:18]
    end
    if (reset) begin // @[ListBuffer.scala 50:22]
      valid <= 4'h0; // @[ListBuffer.scala 50:22]
    end else begin
      valid <= _valid_T_4;
    end
    if (reset) begin // @[ListBuffer.scala 53:22]
      used <= 4'h0; // @[ListBuffer.scala 53:22]
    end else begin
      used <= _used_T_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(~io_pop_valid | _T_4[0])) begin
          $fatal; // @[ListBuffer.scala 101:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_pop_valid | _T_4[0])) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ListBuffer.scala:101 assert (!io.pop.fire() || (io.valid)(io.pop.bits))\n"); // @[ListBuffer.scala 101:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8 & ~(~io_pop2_valid | _T_11[0])) begin
          $fatal; // @[ListBuffer.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~io_pop2_valid | _T_11[0])) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ListBuffer.scala:103 assert(!io.pop2.get.fire()||(io.valid)(io.pop2.get.bits))\n"
            ); // @[ListBuffer.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    head[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    tail[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    next[initvar] = _RAND_2[1:0];
  _RAND_3 = {9{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data[initvar] = _RAND_3[263:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  valid = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  used = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkA(
  input          clock,
  input          reset,
  input          io_req_ready,
  output         io_req_valid,
  output [2:0]   io_req_bits_opcode,
  output [3:0]   io_req_bits_source,
  output [25:0]  io_req_bits_tag,
  output [4:0]   io_req_bits_offset,
  output [1:0]   io_req_bits_put,
  output [255:0] io_req_bits_data,
  output [7:0]   io_req_bits_mask,
  output         io_req_bits_set,
  output         io_a_ready,
  input          io_a_valid,
  input  [2:0]   io_a_bits_opcode,
  input  [3:0]   io_a_bits_source,
  input  [31:0]  io_a_bits_address,
  input  [31:0]  io_a_bits_mask,
  input  [255:0] io_a_bits_data,
  output         io_pb_pop_ready,
  input          io_pb_pop_valid,
  input  [1:0]   io_pb_pop_bits_index,
  output [255:0] io_pb_beat_data,
  output [7:0]   io_pb_beat_mask,
  output         io_pb_pop2_ready,
  input          io_pb_pop2_valid,
  input  [1:0]   io_pb_pop2_bits_index,
  output [255:0] io_pb_beat2_data,
  output [7:0]   io_pb_beat2_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  putbuffer_clock; // @[SinkA.scala 54:25]
  wire  putbuffer_reset; // @[SinkA.scala 54:25]
  wire  putbuffer_io_push_ready; // @[SinkA.scala 54:25]
  wire  putbuffer_io_push_valid; // @[SinkA.scala 54:25]
  wire [1:0] putbuffer_io_push_bits_index; // @[SinkA.scala 54:25]
  wire [255:0] putbuffer_io_push_bits_data_data; // @[SinkA.scala 54:25]
  wire [7:0] putbuffer_io_push_bits_data_mask; // @[SinkA.scala 54:25]
  wire [3:0] putbuffer_io_valid; // @[SinkA.scala 54:25]
  wire  putbuffer_io_pop_valid; // @[SinkA.scala 54:25]
  wire [1:0] putbuffer_io_pop_bits; // @[SinkA.scala 54:25]
  wire [255:0] putbuffer_io_data_data; // @[SinkA.scala 54:25]
  wire [7:0] putbuffer_io_data_mask; // @[SinkA.scala 54:25]
  wire  putbuffer_io_pop2_valid; // @[SinkA.scala 54:25]
  wire [1:0] putbuffer_io_pop2_bits; // @[SinkA.scala 54:25]
  wire [255:0] putbuffer_io_data2_data; // @[SinkA.scala 54:25]
  wire [7:0] putbuffer_io_data2_mask; // @[SinkA.scala 54:25]
  reg [3:0] lists; // @[SinkA.scala 55:22]
  wire  hasData = io_a_bits_opcode == 3'h0 | io_a_bits_opcode == 3'h1; // @[Parameters.scala 168:23]
  wire  req_block = ~io_req_ready; // @[SinkA.scala 72:19]
  wire  _T_1 = ~req_block; // @[SinkA.scala 80:31]
  wire  _T_2 = io_a_valid & hasData & ~req_block; // @[SinkA.scala 80:28]
  wire  buf_block = hasData & ~putbuffer_io_push_ready; // @[SinkA.scala 73:27]
  wire  _T_3 = ~buf_block; // @[SinkA.scala 80:45]
  wire [3:0] _freeOH_T = ~lists; // @[SinkA.scala 63:23]
  wire [4:0] _freeOH_T_1 = {_freeOH_T, 1'h0}; // @[package.scala 244:48]
  wire [3:0] _freeOH_T_3 = _freeOH_T | _freeOH_T_1[3:0]; // @[package.scala 244:43]
  wire [5:0] _freeOH_T_4 = {_freeOH_T_3, 2'h0}; // @[package.scala 244:48]
  wire [3:0] _freeOH_T_6 = _freeOH_T_3 | _freeOH_T_4[3:0]; // @[package.scala 244:43]
  wire [4:0] _freeOH_T_8 = {_freeOH_T_6, 1'h0}; // @[SinkA.scala 63:41]
  wire [4:0] _freeOH_T_9 = ~_freeOH_T_8; // @[SinkA.scala 63:13]
  wire [4:0] _GEN_4 = {{1'd0}, _freeOH_T}; // @[SinkA.scala 63:57]
  wire [4:0] _freeOH_T_11 = _freeOH_T_9 & _GEN_4; // @[SinkA.scala 63:57]
  wire [3:0] freeOH = _freeOH_T_11[3:0]; // @[SinkA.scala 62:20 63:10]
  wire [3:0] lists_set = io_a_valid & hasData & ~req_block & ~buf_block ? freeOH : 4'h0; // @[SinkA.scala 80:{57,69}]
  wire [3:0] _lists_T = lists | lists_set; // @[SinkA.scala 59:19]
  wire  _T_5 = io_pb_pop_ready & io_pb_pop_valid; // @[Decoupled.scala 50:35]
  wire  _T_6 = io_pb_pop2_ready & io_pb_pop2_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _lists_clr_T = 4'h1 << io_pb_pop_bits_index; // @[OneHot.scala 64:12]
  wire [3:0] _lists_clr_T_2 = 4'h1 << io_pb_pop2_bits_index; // @[OneHot.scala 64:12]
  wire [3:0] _lists_clr_T_4 = _lists_clr_T | _lists_clr_T_2; // @[SinkA.scala 110:70]
  wire [3:0] _GEN_1 = _T_6 ? _lists_clr_T_4 : _lists_clr_T; // @[SinkA.scala 109:30 110:19 111:19]
  wire [3:0] _GEN_2 = _T_5 ? _GEN_1 : _lists_clr_T_2; // @[SinkA.scala 108:27 113:16]
  wire [3:0] lists_clr = _T_5 | _T_6 ? _GEN_2 : 4'h0; // @[SinkA.scala 107:46]
  wire [3:0] _lists_T_1 = ~lists_clr; // @[SinkA.scala 59:35]
  wire [3:0] _lists_T_2 = _lists_T & _lists_T_1; // @[SinkA.scala 59:32]
  wire  free = ~(&lists); // @[SinkA.scala 61:14]
  wire [1:0] freeIdx_hi = freeOH[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] freeIdx_lo = freeOH[1:0]; // @[OneHot.scala 31:18]
  wire  _freeIdx_T = |freeIdx_hi; // @[OneHot.scala 32:14]
  wire [1:0] _freeIdx_T_1 = freeIdx_hi | freeIdx_lo; // @[OneHot.scala 32:28]
  wire  set_block = hasData & ~free; // @[SinkA.scala 74:27]
  wire  _io_a_ready_T_3 = ~set_block; // @[SinkA.scala 77:42]
  wire [26:0] set = io_a_bits_address[31:5]; // @[Parameters.scala 214:22]
  wire [3:0] _io_pb_pop_ready_T = putbuffer_io_valid >> io_pb_pop_bits_index; // @[SinkA.scala 102:40]
  wire [3:0] _io_pb_pop2_ready_T = putbuffer_io_valid >> io_pb_pop2_bits_index; // @[SinkA.scala 103:40]
  ListBuffer putbuffer ( // @[SinkA.scala 54:25]
    .clock(putbuffer_clock),
    .reset(putbuffer_reset),
    .io_push_ready(putbuffer_io_push_ready),
    .io_push_valid(putbuffer_io_push_valid),
    .io_push_bits_index(putbuffer_io_push_bits_index),
    .io_push_bits_data_data(putbuffer_io_push_bits_data_data),
    .io_push_bits_data_mask(putbuffer_io_push_bits_data_mask),
    .io_valid(putbuffer_io_valid),
    .io_pop_valid(putbuffer_io_pop_valid),
    .io_pop_bits(putbuffer_io_pop_bits),
    .io_data_data(putbuffer_io_data_data),
    .io_data_mask(putbuffer_io_data_mask),
    .io_pop2_valid(putbuffer_io_pop2_valid),
    .io_pop2_bits(putbuffer_io_pop2_bits),
    .io_data2_data(putbuffer_io_data2_data),
    .io_data2_mask(putbuffer_io_data2_mask)
  );
  assign io_req_valid = io_a_valid & _T_3 & _io_a_ready_T_3; // @[SinkA.scala 78:41]
  assign io_req_bits_opcode = io_a_bits_opcode; // @[SinkA.scala 85:22]
  assign io_req_bits_source = io_a_bits_source; // @[SinkA.scala 87:22]
  assign io_req_bits_tag = set[26:1]; // @[Parameters.scala 215:19]
  assign io_req_bits_offset = io_a_bits_address[4:0]; // @[Parameters.scala 216:50]
  assign io_req_bits_put = {_freeIdx_T,_freeIdx_T_1[1]}; // @[Cat.scala 31:58]
  assign io_req_bits_data = io_a_bits_data; // @[SinkA.scala 93:22]
  assign io_req_bits_mask = io_a_bits_mask[7:0]; // @[SinkA.scala 92:22]
  assign io_req_bits_set = set[0]; // @[Parameters.scala 216:28]
  assign io_a_ready = _T_1 & _T_3 & ~set_block; // @[SinkA.scala 77:39]
  assign io_pb_pop_ready = _io_pb_pop_ready_T[0]; // @[SinkA.scala 102:40]
  assign io_pb_beat_data = putbuffer_io_data_data; // @[SinkA.scala 104:14]
  assign io_pb_beat_mask = putbuffer_io_data_mask; // @[SinkA.scala 104:14]
  assign io_pb_pop2_ready = _io_pb_pop2_ready_T[0]; // @[SinkA.scala 103:40]
  assign io_pb_beat2_data = putbuffer_io_data2_data; // @[SinkA.scala 105:14]
  assign io_pb_beat2_mask = putbuffer_io_data2_mask; // @[SinkA.scala 105:14]
  assign putbuffer_clock = clock;
  assign putbuffer_reset = reset;
  assign putbuffer_io_push_valid = _T_2 & _io_a_ready_T_3; // @[SinkA.scala 79:63]
  assign putbuffer_io_push_bits_index = {_freeIdx_T,_freeIdx_T_1[1]}; // @[Cat.scala 31:58]
  assign putbuffer_io_push_bits_data_data = io_a_bits_data; // @[SinkA.scala 95:36]
  assign putbuffer_io_push_bits_data_mask = io_a_bits_mask[7:0]; // @[SinkA.scala 96:36]
  assign putbuffer_io_pop_valid = io_pb_pop_ready & io_pb_pop_valid; // @[Decoupled.scala 50:35]
  assign putbuffer_io_pop_bits = io_pb_pop_bits_index; // @[SinkA.scala 98:25]
  assign putbuffer_io_pop2_valid = io_pb_pop2_ready & io_pb_pop2_valid; // @[Decoupled.scala 50:35]
  assign putbuffer_io_pop2_bits = io_pb_pop2_bits_index; // @[SinkA.scala 100:29]
  always @(posedge clock) begin
    if (reset) begin // @[SinkA.scala 55:22]
      lists <= 4'h0; // @[SinkA.scala 55:22]
    end else begin
      lists <= _lists_T_2; // @[SinkA.scala 59:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lists = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_105(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [2:0]   io_enq_bits_opcode,
  input  [3:0]   io_enq_bits_source,
  input  [255:0] io_enq_bits_data,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [3:0]   io_deq_bits_source,
  output [255:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [255:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [255:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [255:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [255:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      value <= value + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (io_deq_valid) begin // @[Decoupled.scala 276:16]
      value_1 <= value_1 + 1'h1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != io_deq_valid) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_1[3:0];
  _RAND_2 = {8{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[255:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinkD(
  input          clock,
  input          reset,
  output         io_resp_valid,
  output [2:0]   io_resp_bits_opcode,
  output [3:0]   io_resp_bits_source,
  output [255:0] io_resp_bits_data,
  output         io_d_ready,
  input          io_d_valid,
  input  [2:0]   io_d_bits_opcode,
  input  [3:0]   io_d_bits_source,
  input  [255:0] io_d_bits_data,
  output [3:0]   io_source,
  input  [1:0]   io_way,
  input          io_set,
  input  [2:0]   io_opcode,
  input  [1:0]   io_put,
  output         io_bs_adr_valid,
  output [1:0]   io_bs_adr_bits_way,
  output         io_bs_adr_bits_set,
  output [255:0] io_bs_dat_data,
  output         io_pb_pop_valid,
  output [1:0]   io_pb_pop_bits_index,
  input  [255:0] io_pb_beat_data,
  input  [7:0]   io_pb_beat_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  d_clock; // @[Decoupled.scala 361:21]
  wire  d_reset; // @[Decoupled.scala 361:21]
  wire  d_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  d_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] d_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] d_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [255:0] d_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  d_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  d_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] d_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] d_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [255:0] d_io_deq_bits_data; // @[Decoupled.scala 361:21]
  reg [3:0] io_source_r; // @[Reg.scala 16:16]
  wire [31:0] _full_mask_T_9 = io_pb_beat_mask[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_11 = io_pb_beat_mask[1] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_13 = io_pb_beat_mask[2] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_15 = io_pb_beat_mask[3] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_17 = io_pb_beat_mask[4] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_19 = io_pb_beat_mask[5] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_21 = io_pb_beat_mask[6] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _full_mask_T_23 = io_pb_beat_mask[7] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [255:0] full_mask = {_full_mask_T_23,_full_mask_T_21,_full_mask_T_19,_full_mask_T_17,_full_mask_T_15,
    _full_mask_T_13,_full_mask_T_11,_full_mask_T_9}; // @[Cat.scala 31:58]
  wire [255:0] _merge_data_T = io_pb_beat_data & full_mask; // @[SinkD.scala 58:36]
  wire [255:0] _merge_data_T_1 = ~full_mask; // @[SinkD.scala 58:66]
  wire [255:0] _merge_data_T_2 = d_io_deq_bits_data & _merge_data_T_1; // @[SinkD.scala 58:63]
  wire [255:0] merge_data = _merge_data_T | _merge_data_T_2; // @[SinkD.scala 58:49]
  wire  _io_resp_bits_data_T = io_opcode == 3'h1; // @[SinkD.scala 65:40]
  Queue_105 d ( // @[Decoupled.scala 361:21]
    .clock(d_clock),
    .reset(d_reset),
    .io_enq_ready(d_io_enq_ready),
    .io_enq_valid(d_io_enq_valid),
    .io_enq_bits_opcode(d_io_enq_bits_opcode),
    .io_enq_bits_source(d_io_enq_bits_source),
    .io_enq_bits_data(d_io_enq_bits_data),
    .io_deq_ready(d_io_deq_ready),
    .io_deq_valid(d_io_deq_valid),
    .io_deq_bits_opcode(d_io_deq_bits_opcode),
    .io_deq_bits_source(d_io_deq_bits_source),
    .io_deq_bits_data(d_io_deq_bits_data)
  );
  assign io_resp_valid = d_io_deq_ready & d_io_deq_valid; // @[Decoupled.scala 50:35]
  assign io_resp_bits_opcode = d_io_deq_bits_opcode; // @[SinkD.scala 63:23]
  assign io_resp_bits_source = d_io_deq_bits_source; // @[SinkD.scala 64:23]
  assign io_resp_bits_data = io_opcode == 3'h1 ? merge_data : d_io_deq_bits_data; // @[SinkD.scala 65:29]
  assign io_d_ready = d_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_source = d_io_deq_valid ? d_io_deq_bits_source : io_source_r; // @[SinkD.scala 56:19]
  assign io_bs_adr_valid = d_io_deq_valid; // @[SinkD.scala 67:23]
  assign io_bs_adr_bits_way = io_way; // @[SinkD.scala 68:23]
  assign io_bs_adr_bits_set = io_set; // @[SinkD.scala 69:23]
  assign io_bs_dat_data = _io_resp_bits_data_T ? merge_data : d_io_deq_bits_data; // @[SinkD.scala 70:29]
  assign io_pb_pop_valid = (_io_resp_bits_data_T | io_opcode == 3'h0) & d_io_deq_valid; // @[SinkD.scala 72:85]
  assign io_pb_pop_bits_index = io_put; // @[SinkD.scala 73:23]
  assign d_clock = clock;
  assign d_reset = reset;
  assign d_io_enq_valid = io_d_valid; // @[Decoupled.scala 363:22]
  assign d_io_enq_bits_opcode = io_d_bits_opcode; // @[Decoupled.scala 364:21]
  assign d_io_enq_bits_source = io_d_bits_source; // @[Decoupled.scala 364:21]
  assign d_io_enq_bits_data = io_d_bits_data; // @[Decoupled.scala 364:21]
  assign d_io_deq_ready = 1'h1; // @[SinkD.scala 61:23]
  always @(posedge clock) begin
    if (d_io_deq_valid) begin // @[Reg.scala 17:18]
      io_source_r <= d_io_deq_bits_source; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_source_r = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_38(
  input         clock,
  input         reset,
  input         io_r_req_valid,
  input         io_r_req_bits_setIdx,
  output [26:0] io_r_resp_data_0,
  output [26:0] io_r_resp_data_1,
  output [26:0] io_r_resp_data_2,
  output [26:0] io_r_resp_data_3,
  input         io_w_req_valid,
  input         io_w_req_bits_setIdx,
  input  [26:0] io_w_req_bits_data_0,
  input  [26:0] io_w_req_bits_data_1,
  input  [26:0] io_w_req_bits_data_2,
  input  [26:0] io_w_req_bits_data_3,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [26:0] array_0 [0:1]; // @[SRAMTemplate.scala 102:26]
  wire  array_0_raw_rdata_en; // @[SRAMTemplate.scala 102:26]
  wire  array_0_raw_rdata_addr; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_0_raw_rdata_data; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_0_MPORT_data; // @[SRAMTemplate.scala 102:26]
  wire  array_0_MPORT_addr; // @[SRAMTemplate.scala 102:26]
  wire  array_0_MPORT_mask; // @[SRAMTemplate.scala 102:26]
  wire  array_0_MPORT_en; // @[SRAMTemplate.scala 102:26]
  reg  array_0_raw_rdata_en_pipe_0;
  reg  array_0_raw_rdata_addr_pipe_0;
  reg [26:0] array_1 [0:1]; // @[SRAMTemplate.scala 102:26]
  wire  array_1_raw_rdata_en; // @[SRAMTemplate.scala 102:26]
  wire  array_1_raw_rdata_addr; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_1_raw_rdata_data; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_1_MPORT_data; // @[SRAMTemplate.scala 102:26]
  wire  array_1_MPORT_addr; // @[SRAMTemplate.scala 102:26]
  wire  array_1_MPORT_mask; // @[SRAMTemplate.scala 102:26]
  wire  array_1_MPORT_en; // @[SRAMTemplate.scala 102:26]
  reg  array_1_raw_rdata_en_pipe_0;
  reg  array_1_raw_rdata_addr_pipe_0;
  reg [26:0] array_2 [0:1]; // @[SRAMTemplate.scala 102:26]
  wire  array_2_raw_rdata_en; // @[SRAMTemplate.scala 102:26]
  wire  array_2_raw_rdata_addr; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_2_raw_rdata_data; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_2_MPORT_data; // @[SRAMTemplate.scala 102:26]
  wire  array_2_MPORT_addr; // @[SRAMTemplate.scala 102:26]
  wire  array_2_MPORT_mask; // @[SRAMTemplate.scala 102:26]
  wire  array_2_MPORT_en; // @[SRAMTemplate.scala 102:26]
  reg  array_2_raw_rdata_en_pipe_0;
  reg  array_2_raw_rdata_addr_pipe_0;
  reg [26:0] array_3 [0:1]; // @[SRAMTemplate.scala 102:26]
  wire  array_3_raw_rdata_en; // @[SRAMTemplate.scala 102:26]
  wire  array_3_raw_rdata_addr; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_3_raw_rdata_data; // @[SRAMTemplate.scala 102:26]
  wire [26:0] array_3_MPORT_data; // @[SRAMTemplate.scala 102:26]
  wire  array_3_MPORT_addr; // @[SRAMTemplate.scala 102:26]
  wire  array_3_MPORT_mask; // @[SRAMTemplate.scala 102:26]
  wire  array_3_MPORT_en; // @[SRAMTemplate.scala 102:26]
  reg  array_3_raw_rdata_en_pipe_0;
  reg  array_3_raw_rdata_addr_pipe_0;
  reg  resetState; // @[SRAMTemplate.scala 106:30]
  reg  wrap_wrap; // @[Counter.scala 62:40]
  wire  resetFinish = resetState & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[SRAMTemplate.scala 108:24 106:30 108:38]
  wire [3:0] waymask = resetState ? 4'hf : io_w_req_bits_waymask; // @[SRAMTemplate.scala 119:20]
  reg [26:0] bypass_wdata_REG_0; // @[SRAMTemplate.scala 134:54]
  reg [26:0] bypass_wdata_REG_1; // @[SRAMTemplate.scala 134:54]
  reg [26:0] bypass_wdata_REG_2; // @[SRAMTemplate.scala 134:54]
  reg [26:0] bypass_wdata_REG_3; // @[SRAMTemplate.scala 134:54]
  reg  bypass_mask_need_check; // @[SRAMTemplate.scala 127:29]
  reg  bypass_mask_waddr_reg; // @[SRAMTemplate.scala 128:28]
  reg  bypass_mask_raddr_reg; // @[SRAMTemplate.scala 129:28]
  wire  _bypass_mask_bypass_T_1 = bypass_mask_need_check & bypass_mask_waddr_reg == bypass_mask_raddr_reg; // @[SRAMTemplate.scala 131:39]
  wire [3:0] _bypass_mask_bypass_T_3 = _bypass_mask_bypass_T_1 ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  reg [3:0] bypass_mask_bypass_REG; // @[SRAMTemplate.scala 131:76]
  wire [3:0] bypass_mask_bypass = _bypass_mask_bypass_T_3 & bypass_mask_bypass_REG; // @[SRAMTemplate.scala 131:67]
  assign array_0_raw_rdata_en = array_0_raw_rdata_en_pipe_0;
  assign array_0_raw_rdata_addr = array_0_raw_rdata_addr_pipe_0;
  assign array_0_raw_rdata_data = array_0[array_0_raw_rdata_addr]; // @[SRAMTemplate.scala 102:26]
  assign array_0_MPORT_data = resetState ? 27'h0 : io_w_req_bits_data_0;
  assign array_0_MPORT_addr = resetState ? wrap_wrap : io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = waymask[0];
  assign array_0_MPORT_en = io_w_req_valid | resetState;
  assign array_1_raw_rdata_en = array_1_raw_rdata_en_pipe_0;
  assign array_1_raw_rdata_addr = array_1_raw_rdata_addr_pipe_0;
  assign array_1_raw_rdata_data = array_1[array_1_raw_rdata_addr]; // @[SRAMTemplate.scala 102:26]
  assign array_1_MPORT_data = resetState ? 27'h0 : io_w_req_bits_data_1;
  assign array_1_MPORT_addr = resetState ? wrap_wrap : io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = waymask[1];
  assign array_1_MPORT_en = io_w_req_valid | resetState;
  assign array_2_raw_rdata_en = array_2_raw_rdata_en_pipe_0;
  assign array_2_raw_rdata_addr = array_2_raw_rdata_addr_pipe_0;
  assign array_2_raw_rdata_data = array_2[array_2_raw_rdata_addr]; // @[SRAMTemplate.scala 102:26]
  assign array_2_MPORT_data = resetState ? 27'h0 : io_w_req_bits_data_2;
  assign array_2_MPORT_addr = resetState ? wrap_wrap : io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = waymask[2];
  assign array_2_MPORT_en = io_w_req_valid | resetState;
  assign array_3_raw_rdata_en = array_3_raw_rdata_en_pipe_0;
  assign array_3_raw_rdata_addr = array_3_raw_rdata_addr_pipe_0;
  assign array_3_raw_rdata_data = array_3[array_3_raw_rdata_addr]; // @[SRAMTemplate.scala 102:26]
  assign array_3_MPORT_data = resetState ? 27'h0 : io_w_req_bits_data_3;
  assign array_3_MPORT_addr = resetState ? wrap_wrap : io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = waymask[3];
  assign array_3_MPORT_en = io_w_req_valid | resetState;
  assign io_r_resp_data_0 = bypass_mask_bypass[0] ? bypass_wdata_REG_0 : array_0_raw_rdata_data; // @[SRAMTemplate.scala 140:30]
  assign io_r_resp_data_1 = bypass_mask_bypass[1] ? bypass_wdata_REG_1 : array_1_raw_rdata_data; // @[SRAMTemplate.scala 140:30]
  assign io_r_resp_data_2 = bypass_mask_bypass[2] ? bypass_wdata_REG_2 : array_2_raw_rdata_data; // @[SRAMTemplate.scala 140:30]
  assign io_r_resp_data_3 = bypass_mask_bypass[3] ? bypass_wdata_REG_3 : array_3_raw_rdata_data; // @[SRAMTemplate.scala 140:30]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[SRAMTemplate.scala 102:26]
    end
    array_0_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_0_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[SRAMTemplate.scala 102:26]
    end
    array_1_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_1_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[SRAMTemplate.scala 102:26]
    end
    array_2_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_2_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[SRAMTemplate.scala 102:26]
    end
    array_3_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_3_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2; // @[SRAMTemplate.scala 106:{30,30}]
    if (reset) begin // @[Counter.scala 62:40]
      wrap_wrap <= 1'h0; // @[Counter.scala 62:40]
    end else if (resetState) begin // @[Counter.scala 120:16]
      wrap_wrap <= wrap_wrap + 1'h1; // @[Counter.scala 78:15]
    end
    bypass_wdata_REG_0 <= io_w_req_bits_data_0; // @[SRAMTemplate.scala 134:54]
    bypass_wdata_REG_1 <= io_w_req_bits_data_1; // @[SRAMTemplate.scala 134:54]
    bypass_wdata_REG_2 <= io_w_req_bits_data_2; // @[SRAMTemplate.scala 134:54]
    bypass_wdata_REG_3 <= io_w_req_bits_data_3; // @[SRAMTemplate.scala 134:54]
    bypass_mask_need_check <= io_r_req_valid & io_w_req_valid; // @[SRAMTemplate.scala 127:34]
    bypass_mask_waddr_reg <= io_w_req_bits_setIdx; // @[SRAMTemplate.scala 128:28]
    bypass_mask_raddr_reg <= io_r_req_bits_setIdx; // @[SRAMTemplate.scala 129:28]
    bypass_mask_bypass_REG <= io_w_req_bits_waymask; // @[SRAMTemplate.scala 131:76]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    array_0[initvar] = _RAND_0[26:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    array_1[initvar] = _RAND_3[26:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    array_2[initvar] = _RAND_6[26:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    array_3[initvar] = _RAND_9[26:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_raw_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_raw_rdata_addr_pipe_0 = _RAND_2[0:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_raw_rdata_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_raw_rdata_addr_pipe_0 = _RAND_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_raw_rdata_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_raw_rdata_addr_pipe_0 = _RAND_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_raw_rdata_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_raw_rdata_addr_pipe_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  resetState = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  wrap_wrap = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bypass_wdata_REG_0 = _RAND_14[26:0];
  _RAND_15 = {1{`RANDOM}};
  bypass_wdata_REG_1 = _RAND_15[26:0];
  _RAND_16 = {1{`RANDOM}};
  bypass_wdata_REG_2 = _RAND_16[26:0];
  _RAND_17 = {1{`RANDOM}};
  bypass_wdata_REG_3 = _RAND_17[26:0];
  _RAND_18 = {1{`RANDOM}};
  bypass_mask_need_check = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  bypass_mask_waddr_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  bypass_mask_raddr_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  bypass_mask_bypass_REG = _RAND_21[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Directory_test(
  input          clock,
  input          reset,
  output         io_write_ready,
  input          io_write_valid,
  input  [1:0]   io_write_bits_way,
  input  [25:0]  io_write_bits_data_tag,
  input          io_write_bits_data_valid,
  input          io_write_bits_set,
  output         io_read_ready,
  input          io_read_valid,
  input  [2:0]   io_read_bits_opcode,
  input  [3:0]   io_read_bits_source,
  input  [25:0]  io_read_bits_tag,
  input  [4:0]   io_read_bits_offset,
  input  [1:0]   io_read_bits_put,
  input  [255:0] io_read_bits_data,
  input  [7:0]   io_read_bits_mask,
  input          io_read_bits_set,
  output         io_result_valid,
  output [2:0]   io_result_bits_opcode,
  output [3:0]   io_result_bits_source,
  output [25:0]  io_result_bits_tag,
  output [4:0]   io_result_bits_offset,
  output [1:0]   io_result_bits_put,
  output [255:0] io_result_bits_data,
  output [7:0]   io_result_bits_mask,
  output         io_result_bits_set,
  output         io_result_bits_hit,
  output [1:0]   io_result_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [255:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  cc_dir_clock; // @[Directory_test.scala 73:22]
  wire  cc_dir_reset; // @[Directory_test.scala 73:22]
  wire  cc_dir_io_r_req_valid; // @[Directory_test.scala 73:22]
  wire  cc_dir_io_r_req_bits_setIdx; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_r_resp_data_0; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_r_resp_data_1; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_r_resp_data_2; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_r_resp_data_3; // @[Directory_test.scala 73:22]
  wire  cc_dir_io_w_req_valid; // @[Directory_test.scala 73:22]
  wire  cc_dir_io_w_req_bits_setIdx; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_w_req_bits_data_0; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_w_req_bits_data_1; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_w_req_bits_data_2; // @[Directory_test.scala 73:22]
  wire [26:0] cc_dir_io_w_req_bits_data_3; // @[Directory_test.scala 73:22]
  wire [3:0] cc_dir_io_w_req_bits_waymask; // @[Directory_test.scala 73:22]
  reg [1:0] wipeCount; // @[Directory_test.scala 81:26]
  reg  wipeOff; // @[Directory_test.scala 82:26]
  wire  wipeDone = wipeCount[1]; // @[Directory_test.scala 83:28]
  wire  wipeSet = wipeCount[0]; // @[Directory_test.scala 84:28]
  wire  _T = ~wipeDone; // @[Directory_test.scala 89:9]
  wire  _T_2 = ~wipeDone & ~wipeOff; // @[Directory_test.scala 89:19]
  wire [1:0] _wipeCount_T_1 = wipeCount + 2'h1; // @[Directory_test.scala 89:57]
  wire  ren = io_read_ready & io_read_valid; // @[Decoupled.scala 50:35]
  wire  _wen_new_T_3 = io_write_ready & io_write_valid; // @[Decoupled.scala 50:35]
  reg  ren1; // @[Directory_test.scala 102:21]
  reg  wen1; // @[Directory_test.scala 104:19]
  reg [25:0] tag; // @[Reg.scala 16:16]
  reg  set; // @[Reg.scala 16:16]
  reg  state_reg; // @[Replacement.scala 168:70]
  reg  state_reg_1; // @[Replacement.scala 168:70]
  wire  setQuash_1 = _wen_new_T_3 & io_write_bits_set == io_read_bits_set; // @[Directory_test.scala 120:24]
  wire  setQuash = wen1 & io_write_bits_set == set; // @[Directory_test.scala 121:21]
  wire  tagMatch_1 = io_write_bits_data_tag == io_read_bits_tag; // @[Directory_test.scala 122:41]
  wire  tagMatch = io_write_bits_data_tag == tag; // @[Directory_test.scala 123:41]
  reg [1:0] writeWay1; // @[Directory_test.scala 124:26]
  wire [107:0] _ways_T = {cc_dir_io_r_resp_data_3,cc_dir_io_r_resp_data_2,cc_dir_io_r_resp_data_1,
    cc_dir_io_r_resp_data_0}; // @[Directory_test.scala 126:29]
  wire  ways_0_valid = _ways_T[0]; // @[Directory_test.scala 126:29]
  wire [25:0] ways_0_tag = _ways_T[26:1]; // @[Directory_test.scala 126:29]
  wire  ways_1_valid = _ways_T[27]; // @[Directory_test.scala 126:29]
  wire [25:0] ways_1_tag = _ways_T[53:28]; // @[Directory_test.scala 126:29]
  wire  ways_2_valid = _ways_T[54]; // @[Directory_test.scala 126:29]
  wire [25:0] ways_2_tag = _ways_T[80:55]; // @[Directory_test.scala 126:29]
  wire  ways_3_valid = _ways_T[81]; // @[Directory_test.scala 126:29]
  wire [25:0] ways_3_tag = _ways_T[107:82]; // @[Directory_test.scala 126:29]
  wire  _hits_T_3 = ways_0_tag == tag & ~setQuash & ways_0_valid; // @[Directory_test.scala 129:35]
  wire  _hits_T_7 = ways_1_tag == tag & ~setQuash & ways_1_valid; // @[Directory_test.scala 129:35]
  wire  _hits_T_11 = ways_2_tag == tag & ~setQuash & ways_2_valid; // @[Directory_test.scala 129:35]
  wire  _hits_T_15 = ways_3_tag == tag & ~setQuash & ways_3_valid; // @[Directory_test.scala 129:35]
  wire [3:0] hits = {_hits_T_15,_hits_T_11,_hits_T_7,_hits_T_3}; // @[Cat.scala 31:58]
  wire  _cc_dir_io_r_req_valid_T = setQuash_1 & tagMatch_1; // @[Directory_test.scala 139:48]
  wire  hit = |hits; // @[Directory_test.scala 144:21]
  wire [1:0] hitWay_hi = hits[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] hitWay_lo = hits[1:0]; // @[OneHot.scala 31:18]
  wire  _hitWay_T = |hitWay_hi; // @[OneHot.scala 32:14]
  wire [1:0] _hitWay_T_1 = hitWay_hi | hitWay_lo; // @[OneHot.scala 32:28]
  wire [1:0] hitWay = {_hitWay_T,_hitWay_T_1[1]}; // @[Cat.scala 31:58]
  reg  writeSet1; // @[Directory_test.scala 147:26]
  wire  state_reg_touch_way_sized = writeWay1[0]; // @[package.scala 154:13]
  wire  _state_reg_T_1 = ~state_reg_touch_way_sized; // @[Replacement.scala 218:7]
  wire  state_reg_touch_way_sized_1 = hitWay[0]; // @[package.scala 154:13]
  wire  _state_reg_T_3 = ~state_reg_touch_way_sized_1; // @[Replacement.scala 218:7]
  wire [26:0] _x5_T = {io_write_bits_data_tag,io_write_bits_data_valid}; // @[Directory_test.scala 161:43]
  wire  x6_shiftAmount = io_write_bits_way[0]; // @[OneHot.scala 63:49]
  wire [1:0] _x6_T = 2'h1 << x6_shiftAmount; // @[OneHot.scala 64:12]
  wire [1:0] _x6_T_4 = _T ? 2'h3 : 2'h0; // @[Bitwise.scala 74:12]
  wire [1:0] x6 = _x6_T | _x6_T_4; // @[Directory_test.scala 162:44]
  wire  _io_result_bits_hit_T = setQuash & tagMatch; // @[Directory_test.scala 166:42]
  wire  _GEN_8 = set ? state_reg_1 : state_reg; // @[Directory_test.scala 167:{54,54}]
  wire [1:0] _io_result_bits_way_T_5 = _io_result_bits_hit_T ? io_write_bits_way : {{1'd0}, _GEN_8}; // @[Directory_test.scala 167:54]
  reg [1:0] io_result_bits_put_REG; // @[Directory_test.scala 168:34]
  reg [255:0] io_result_bits_data_REG; // @[Directory_test.scala 169:34]
  reg [4:0] io_result_bits_offset_REG; // @[Directory_test.scala 170:34]
  reg  io_result_bits_set_REG; // @[Directory_test.scala 172:34]
  reg [3:0] io_result_bits_source_REG; // @[Directory_test.scala 173:34]
  reg [25:0] io_result_bits_tag_REG; // @[Directory_test.scala 174:34]
  reg [2:0] io_result_bits_opcode_REG; // @[Directory_test.scala 175:34]
  reg [7:0] io_result_bits_mask_REG; // @[Directory_test.scala 176:34]
  SRAMTemplate_38 cc_dir ( // @[Directory_test.scala 73:22]
    .clock(cc_dir_clock),
    .reset(cc_dir_reset),
    .io_r_req_valid(cc_dir_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_dir_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_dir_io_r_resp_data_0),
    .io_r_resp_data_1(cc_dir_io_r_resp_data_1),
    .io_r_resp_data_2(cc_dir_io_r_resp_data_2),
    .io_r_resp_data_3(cc_dir_io_r_resp_data_3),
    .io_w_req_valid(cc_dir_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_dir_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_dir_io_w_req_bits_data_0),
    .io_w_req_bits_data_1(cc_dir_io_w_req_bits_data_1),
    .io_w_req_bits_data_2(cc_dir_io_w_req_bits_data_2),
    .io_w_req_bits_data_3(cc_dir_io_w_req_bits_data_3),
    .io_w_req_bits_waymask(cc_dir_io_w_req_bits_waymask)
  );
  assign io_write_ready = wipeCount[1]; // @[Directory_test.scala 83:28]
  assign io_read_ready = wipeDone & ~_wen_new_T_3 | _cc_dir_io_r_req_valid_T; // @[Directory_test.scala 164:49]
  assign io_result_valid = ren1; // @[Directory_test.scala 165:19]
  assign io_result_bits_opcode = io_result_bits_opcode_REG; // @[Directory_test.scala 175:25]
  assign io_result_bits_source = io_result_bits_source_REG; // @[Directory_test.scala 173:25]
  assign io_result_bits_tag = io_result_bits_tag_REG; // @[Directory_test.scala 174:25]
  assign io_result_bits_offset = io_result_bits_offset_REG; // @[Directory_test.scala 170:25]
  assign io_result_bits_put = io_result_bits_put_REG; // @[Directory_test.scala 168:25]
  assign io_result_bits_data = io_result_bits_data_REG; // @[Directory_test.scala 169:25]
  assign io_result_bits_mask = io_result_bits_mask_REG; // @[Directory_test.scala 176:25]
  assign io_result_bits_set = io_result_bits_set_REG; // @[Directory_test.scala 172:25]
  assign io_result_bits_hit = hit | setQuash & tagMatch; // @[Directory_test.scala 166:30]
  assign io_result_bits_way = hit ? hitWay : _io_result_bits_way_T_5; // @[Directory_test.scala 167:29]
  assign cc_dir_clock = clock;
  assign cc_dir_reset = reset;
  assign cc_dir_io_r_req_valid = ren & ~(setQuash_1 & tagMatch_1); // @[Directory_test.scala 139:32]
  assign cc_dir_io_r_req_bits_setIdx = io_read_bits_set; // @[SRAMTemplate.scala 43:17]
  assign cc_dir_io_w_req_valid = _T_2 | _wen_new_T_3; // @[Directory_test.scala 92:41]
  assign cc_dir_io_w_req_bits_setIdx = wipeDone ? io_write_bits_set : wipeSet; // @[Directory_test.scala 160:15]
  assign cc_dir_io_w_req_bits_data_0 = wipeDone ? _x5_T : 27'h0; // @[Directory_test.scala 161:13]
  assign cc_dir_io_w_req_bits_data_1 = wipeDone ? _x5_T : 27'h0; // @[Directory_test.scala 161:13]
  assign cc_dir_io_w_req_bits_data_2 = wipeDone ? _x5_T : 27'h0; // @[Directory_test.scala 161:13]
  assign cc_dir_io_w_req_bits_data_3 = wipeDone ? _x5_T : 27'h0; // @[Directory_test.scala 161:13]
  assign cc_dir_io_w_req_bits_waymask = {{2'd0}, x6}; // @[SRAMTemplate.scala 55:24]
  always @(posedge clock) begin
    if (reset) begin // @[Directory_test.scala 81:26]
      wipeCount <= 2'h0; // @[Directory_test.scala 81:26]
    end else if (~wipeDone & ~wipeOff) begin // @[Directory_test.scala 89:32]
      wipeCount <= _wipeCount_T_1; // @[Directory_test.scala 89:44]
    end
    wipeOff <= reset; // @[Directory_test.scala 82:{26,26,26}]
    if (reset) begin // @[Directory_test.scala 102:21]
      ren1 <= 1'h0; // @[Directory_test.scala 102:21]
    end else begin
      ren1 <= ren; // @[Directory_test.scala 103:8]
    end
    if (reset) begin // @[Directory_test.scala 104:19]
      wen1 <= 1'h0; // @[Directory_test.scala 104:19]
    end else begin
      wen1 <= _wen_new_T_3; // @[Directory_test.scala 105:7]
    end
    if (ren) begin // @[Reg.scala 17:18]
      tag <= io_read_bits_tag; // @[Reg.scala 17:22]
    end
    if (ren) begin // @[Reg.scala 17:18]
      set <= io_read_bits_set; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Replacement.scala 168:70]
      state_reg <= 1'h0; // @[Replacement.scala 168:70]
    end else if (wen1 & ~writeSet1) begin // @[Directory_test.scala 151:32]
      state_reg <= _state_reg_T_1; // @[Replacement.scala 172:15]
    end else if (ren1 & ~set & hit) begin // @[Directory_test.scala 153:37]
      state_reg <= _state_reg_T_3; // @[Replacement.scala 172:15]
    end
    if (reset) begin // @[Replacement.scala 168:70]
      state_reg_1 <= 1'h0; // @[Replacement.scala 168:70]
    end else if (wen1 & writeSet1) begin // @[Directory_test.scala 151:32]
      state_reg_1 <= _state_reg_T_1; // @[Replacement.scala 172:15]
    end else if (ren1 & set & hit) begin // @[Directory_test.scala 153:37]
      state_reg_1 <= _state_reg_T_3; // @[Replacement.scala 172:15]
    end
    if (reset) begin // @[Directory_test.scala 124:26]
      writeWay1 <= 2'h0; // @[Directory_test.scala 124:26]
    end else begin
      writeWay1 <= io_write_bits_way; // @[Directory_test.scala 125:12]
    end
    writeSet1 <= io_write_bits_set; // @[Directory_test.scala 147:26]
    io_result_bits_put_REG <= io_read_bits_put; // @[Directory_test.scala 168:34]
    io_result_bits_data_REG <= io_read_bits_data; // @[Directory_test.scala 169:34]
    io_result_bits_offset_REG <= io_read_bits_offset; // @[Directory_test.scala 170:34]
    io_result_bits_set_REG <= io_read_bits_set; // @[Directory_test.scala 172:34]
    io_result_bits_source_REG <= io_read_bits_source; // @[Directory_test.scala 173:34]
    io_result_bits_tag_REG <= io_read_bits_tag; // @[Directory_test.scala 174:34]
    io_result_bits_opcode_REG <= io_read_bits_opcode; // @[Directory_test.scala 175:34]
    io_result_bits_mask_REG <= io_read_bits_mask; // @[Directory_test.scala 176:34]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wipeCount = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wipeOff = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ren1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wen1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  tag = _RAND_4[25:0];
  _RAND_5 = {1{`RANDOM}};
  set = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_reg_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  writeWay1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  writeSet1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_result_bits_put_REG = _RAND_10[1:0];
  _RAND_11 = {8{`RANDOM}};
  io_result_bits_data_REG = _RAND_11[255:0];
  _RAND_12 = {1{`RANDOM}};
  io_result_bits_offset_REG = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  io_result_bits_set_REG = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  io_result_bits_source_REG = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  io_result_bits_tag_REG = _RAND_15[25:0];
  _RAND_16 = {1{`RANDOM}};
  io_result_bits_opcode_REG = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  io_result_bits_mask_REG = _RAND_17[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_39(
  input         clock,
  input         reset,
  input         io_r_req_valid,
  input  [1:0]  io_r_req_bits_setIdx,
  output [31:0] io_r_resp_data_0,
  input         io_w_req_valid,
  input  [1:0]  io_w_req_bits_setIdx,
  input  [31:0] io_w_req_bits_data_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] array_0 [0:3]; // @[SRAMTemplate.scala 102:26]
  wire  array_0_raw_rdata_en; // @[SRAMTemplate.scala 102:26]
  wire [1:0] array_0_raw_rdata_addr; // @[SRAMTemplate.scala 102:26]
  wire [31:0] array_0_raw_rdata_data; // @[SRAMTemplate.scala 102:26]
  wire [31:0] array_0_MPORT_data; // @[SRAMTemplate.scala 102:26]
  wire [1:0] array_0_MPORT_addr; // @[SRAMTemplate.scala 102:26]
  wire  array_0_MPORT_mask; // @[SRAMTemplate.scala 102:26]
  wire  array_0_MPORT_en; // @[SRAMTemplate.scala 102:26]
  reg  array_0_raw_rdata_en_pipe_0;
  reg [1:0] array_0_raw_rdata_addr_pipe_0;
  reg  resetState; // @[SRAMTemplate.scala 106:30]
  reg [1:0] resetSet; // @[Counter.scala 62:40]
  wire  wrap_wrap = resetSet == 2'h3; // @[Counter.scala 74:24]
  wire [1:0] _wrap_value_T_1 = resetSet + 2'h1; // @[Counter.scala 78:24]
  wire  resetFinish = resetState & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[SRAMTemplate.scala 108:24 106:30 108:38]
  reg [63:0] bypass_wdata_lfsr; // @[Fuzzer.scala 43:19]
  wire  bypass_wdata_xor = bypass_wdata_lfsr[0] ^ bypass_wdata_lfsr[1] ^ bypass_wdata_lfsr[3] ^ bypass_wdata_lfsr[4]; // @[Fuzzer.scala 44:43]
  wire [63:0] _bypass_wdata_lfsr_T_2 = {bypass_wdata_xor,bypass_wdata_lfsr[63:1]}; // @[Cat.scala 31:58]
  reg  bypass_mask_need_check; // @[SRAMTemplate.scala 127:29]
  reg [1:0] bypass_mask_waddr_reg; // @[SRAMTemplate.scala 128:28]
  reg [1:0] bypass_mask_raddr_reg; // @[SRAMTemplate.scala 129:28]
  wire  bypass_mask_bypass = bypass_mask_need_check & bypass_mask_waddr_reg == bypass_mask_raddr_reg; // @[SRAMTemplate.scala 131:39]
  wire [31:0] bypass_wdata_0 = bypass_wdata_lfsr[31:0]; // @[SRAMTemplate.scala 135:{58,58}]
  assign array_0_raw_rdata_en = array_0_raw_rdata_en_pipe_0;
  assign array_0_raw_rdata_addr = array_0_raw_rdata_addr_pipe_0;
  assign array_0_raw_rdata_data = array_0[array_0_raw_rdata_addr]; // @[SRAMTemplate.scala 102:26]
  assign array_0_MPORT_data = resetState ? 32'h0 : io_w_req_bits_data_0;
  assign array_0_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = 1'h1;
  assign array_0_MPORT_en = io_w_req_valid | resetState;
  assign io_r_resp_data_0 = bypass_mask_bypass ? bypass_wdata_0 : array_0_raw_rdata_data; // @[SRAMTemplate.scala 140:30]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[SRAMTemplate.scala 102:26]
    end
    array_0_raw_rdata_en_pipe_0 <= io_r_req_valid;
    if (io_r_req_valid) begin
      array_0_raw_rdata_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2; // @[SRAMTemplate.scala 106:{30,30}]
    if (reset) begin // @[Counter.scala 62:40]
      resetSet <= 2'h0; // @[Counter.scala 62:40]
    end else if (resetState) begin // @[Counter.scala 120:16]
      resetSet <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
    if (bypass_wdata_lfsr == 64'h0) begin // @[Fuzzer.scala 46:18]
      bypass_wdata_lfsr <= 64'h1;
    end else begin
      bypass_wdata_lfsr <= _bypass_wdata_lfsr_T_2;
    end
    bypass_mask_need_check <= io_r_req_valid & io_w_req_valid; // @[SRAMTemplate.scala 127:34]
    bypass_mask_waddr_reg <= io_w_req_bits_setIdx; // @[SRAMTemplate.scala 128:28]
    bypass_mask_raddr_reg <= io_r_req_bits_setIdx; // @[SRAMTemplate.scala 129:28]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    array_0[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_raw_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_raw_rdata_addr_pipe_0 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  resetState = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  resetSet = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  bypass_wdata_lfsr = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  bypass_mask_need_check = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bypass_mask_waddr_reg = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  bypass_mask_raddr_reg = _RAND_8[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BankedStore(
  input          clock,
  input          reset,
  input          io_sinkD_adr_valid,
  input  [1:0]   io_sinkD_adr_bits_way,
  input          io_sinkD_adr_bits_set,
  input  [255:0] io_sinkD_dat_data,
  input          io_sourceD_radr_valid,
  input  [1:0]   io_sourceD_radr_bits_way,
  input          io_sourceD_radr_bits_set,
  input  [7:0]   io_sourceD_radr_bits_mask,
  output [255:0] io_sourceD_rdat_data,
  input          io_sourceD_wadr_valid,
  input  [1:0]   io_sourceD_wadr_bits_way,
  input          io_sourceD_wadr_bits_set,
  input  [7:0]   io_sourceD_wadr_bits_mask,
  input  [255:0] io_sourceD_wdat_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  cc_banks_0_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_0_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_0_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_0_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_0_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_0_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_0_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_0_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_1_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_1_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_1_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_1_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_1_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_1_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_1_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_1_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_2_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_2_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_2_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_2_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_2_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_2_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_2_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_2_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_3_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_3_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_3_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_3_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_3_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_3_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_3_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_3_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_4_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_4_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_4_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_4_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_4_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_4_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_4_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_4_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_5_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_5_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_5_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_5_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_5_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_5_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_5_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_5_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_6_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_6_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_6_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_6_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_6_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_6_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_6_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_6_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_7_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_7_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_7_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_7_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_7_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_7_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_7_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_7_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_8_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_8_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_8_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_8_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_8_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_8_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_8_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_8_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_9_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_9_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_9_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_9_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_9_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_9_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_9_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_9_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_10_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_10_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_10_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_10_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_10_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_10_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_10_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_10_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_11_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_11_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_11_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_11_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_11_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_11_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_11_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_11_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_12_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_12_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_12_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_12_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_12_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_12_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_12_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_12_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_13_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_13_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_13_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_13_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_13_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_13_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_13_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_13_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_14_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_14_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_14_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_14_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_14_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_14_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_14_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_14_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_15_clock; // @[BankedStore.scala 101:13]
  wire  cc_banks_15_reset; // @[BankedStore.scala 101:13]
  wire  cc_banks_15_io_r_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_15_io_r_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_15_io_r_resp_data_0; // @[BankedStore.scala 101:13]
  wire  cc_banks_15_io_w_req_valid; // @[BankedStore.scala 101:13]
  wire [1:0] cc_banks_15_io_w_req_bits_setIdx; // @[BankedStore.scala 101:13]
  wire [31:0] cc_banks_15_io_w_req_bits_data_0; // @[BankedStore.scala 101:13]
  wire [31:0] sinkD_req_words_0 = io_sinkD_dat_data[31:0]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_1 = io_sinkD_dat_data[63:32]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_2 = io_sinkD_dat_data[95:64]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_3 = io_sinkD_dat_data[127:96]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_4 = io_sinkD_dat_data[159:128]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_5 = io_sinkD_dat_data[191:160]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_6 = io_sinkD_dat_data[223:192]; // @[BankedStore.scala 139:19]
  wire [31:0] sinkD_req_words_7 = io_sinkD_dat_data[255:224]; // @[BankedStore.scala 139:19]
  wire [2:0] sinkD_req_a = {io_sinkD_adr_bits_way,io_sinkD_adr_bits_set}; // @[Cat.scala 31:58]
  wire  sinkD_req_select_shiftAmount = sinkD_req_a[0]; // @[BankedStore.scala 146:28]
  wire [1:0] sinkD_req_select = 2'h1 << sinkD_req_select_shiftAmount; // @[OneHot.scala 64:12]
  wire [1:0] reqs_0_index = sinkD_req_a[2:1]; // @[BankedStore.scala 151:23]
  wire [7:0] _sinkD_req_out_bankSel_T_3 = sinkD_req_select[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _sinkD_req_out_bankSel_T_5 = sinkD_req_select[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [15:0] _sinkD_req_out_bankSel_T_6 = {_sinkD_req_out_bankSel_T_5,_sinkD_req_out_bankSel_T_3}; // @[Cat.scala 31:58]
  wire [15:0] reqs_0_bankSel = io_sinkD_adr_valid ? _sinkD_req_out_bankSel_T_6 : 16'h0; // @[BankedStore.scala 152:24]
  wire [2:0] sourceD_rreq_a = {io_sourceD_radr_bits_way,io_sourceD_radr_bits_set}; // @[Cat.scala 31:58]
  wire  sourceD_rreq_select_shiftAmount = sourceD_rreq_a[0]; // @[BankedStore.scala 146:28]
  wire [1:0] sourceD_rreq_select = 2'h1 << sourceD_rreq_select_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] sourceD_wreq_a = {io_sourceD_wadr_bits_way,io_sourceD_wadr_bits_set}; // @[Cat.scala 31:58]
  wire  sourceD_wreq_select_shiftAmount = sourceD_wreq_a[0]; // @[BankedStore.scala 146:28]
  wire [1:0] sourceD_wreq_select = 2'h1 << sourceD_wreq_select_shiftAmount; // @[OneHot.scala 64:12]
  wire [7:0] _sourceD_wreq_out_bankSel_T_5 = sourceD_wreq_select[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _sourceD_wreq_out_bankSel_T_3 = sourceD_wreq_select[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [15:0] _sourceD_wreq_out_bankSel_T_6 = {_sourceD_wreq_out_bankSel_T_5,_sourceD_wreq_out_bankSel_T_3}; // @[Cat.scala 31:58]
  wire [15:0] _sourceD_wreq_out_bankSel_T_7 = {io_sourceD_wadr_bits_mask,io_sourceD_wadr_bits_mask}; // @[Cat.scala 31:58]
  wire [15:0] _sourceD_wreq_out_bankSel_T_8 = _sourceD_wreq_out_bankSel_T_6 & _sourceD_wreq_out_bankSel_T_7; // @[BankedStore.scala 152:64]
  wire [15:0] reqs_1_bankSel = io_sourceD_wadr_valid ? _sourceD_wreq_out_bankSel_T_8 : 16'h0; // @[BankedStore.scala 152:24]
  wire [15:0] reqs_2_bankSum = reqs_1_bankSel | reqs_0_bankSel; // @[BankedStore.scala 175:17]
  wire [7:0] _sourceD_rreq_ready_T_1 = reqs_2_bankSum[7:0] & io_sourceD_radr_bits_mask; // @[BankedStore.scala 147:96]
  wire  _sourceD_rreq_ready_T_3 = ~(|_sourceD_rreq_ready_T_1); // @[BankedStore.scala 147:58]
  wire [7:0] _sourceD_rreq_ready_T_5 = reqs_2_bankSum[15:8] & io_sourceD_radr_bits_mask; // @[BankedStore.scala 147:96]
  wire  _sourceD_rreq_ready_T_7 = ~(|_sourceD_rreq_ready_T_5); // @[BankedStore.scala 147:58]
  wire [1:0] sourceD_rreq_ready = {_sourceD_rreq_ready_T_7,_sourceD_rreq_ready_T_3}; // @[Cat.scala 31:58]
  wire [1:0] reqs_2_index = sourceD_rreq_a[2:1]; // @[BankedStore.scala 151:23]
  wire [7:0] _sourceD_rreq_out_bankSel_T_3 = sourceD_rreq_select[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _sourceD_rreq_out_bankSel_T_5 = sourceD_rreq_select[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [15:0] _sourceD_rreq_out_bankSel_T_6 = {_sourceD_rreq_out_bankSel_T_5,_sourceD_rreq_out_bankSel_T_3}; // @[Cat.scala 31:58]
  wire [15:0] _sourceD_rreq_out_bankSel_T_7 = {io_sourceD_radr_bits_mask,io_sourceD_radr_bits_mask}; // @[Cat.scala 31:58]
  wire [15:0] _sourceD_rreq_out_bankSel_T_8 = _sourceD_rreq_out_bankSel_T_6 & _sourceD_rreq_out_bankSel_T_7; // @[BankedStore.scala 152:64]
  wire [15:0] reqs_2_bankSel = io_sourceD_radr_valid ? _sourceD_rreq_out_bankSel_T_8 : 16'h0; // @[BankedStore.scala 152:24]
  wire [7:0] _sourceD_rreq_out_bankEn_T_3 = sourceD_rreq_ready[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _sourceD_rreq_out_bankEn_T_5 = sourceD_rreq_ready[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [15:0] _sourceD_rreq_out_bankEn_T_6 = {_sourceD_rreq_out_bankEn_T_5,_sourceD_rreq_out_bankEn_T_3}; // @[Cat.scala 31:58]
  wire [15:0] reqs_2_bankEn = reqs_2_bankSel & _sourceD_rreq_out_bankEn_T_6; // @[BankedStore.scala 153:34]
  wire [31:0] sourceD_wreq_words_0 = io_sourceD_wdat_data[31:0]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_1 = io_sourceD_wdat_data[63:32]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_2 = io_sourceD_wdat_data[95:64]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_3 = io_sourceD_wdat_data[127:96]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_4 = io_sourceD_wdat_data[159:128]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_5 = io_sourceD_wdat_data[191:160]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_6 = io_sourceD_wdat_data[223:192]; // @[BankedStore.scala 139:19]
  wire [31:0] sourceD_wreq_words_7 = io_sourceD_wdat_data[255:224]; // @[BankedStore.scala 139:19]
  wire [7:0] _sourceD_wreq_ready_T_1 = reqs_0_bankSel[7:0] & io_sourceD_wadr_bits_mask; // @[BankedStore.scala 147:96]
  wire  _sourceD_wreq_ready_T_3 = ~(|_sourceD_wreq_ready_T_1); // @[BankedStore.scala 147:58]
  wire [7:0] _sourceD_wreq_ready_T_5 = reqs_0_bankSel[15:8] & io_sourceD_wadr_bits_mask; // @[BankedStore.scala 147:96]
  wire  _sourceD_wreq_ready_T_7 = ~(|_sourceD_wreq_ready_T_5); // @[BankedStore.scala 147:58]
  wire [1:0] sourceD_wreq_ready = {_sourceD_wreq_ready_T_7,_sourceD_wreq_ready_T_3}; // @[Cat.scala 31:58]
  wire [1:0] reqs_1_index = sourceD_wreq_a[2:1]; // @[BankedStore.scala 151:23]
  wire [7:0] _sourceD_wreq_out_bankEn_T_3 = sourceD_wreq_ready[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _sourceD_wreq_out_bankEn_T_5 = sourceD_wreq_ready[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [15:0] _sourceD_wreq_out_bankEn_T_6 = {_sourceD_wreq_out_bankEn_T_5,_sourceD_wreq_out_bankEn_T_3}; // @[Cat.scala 31:58]
  wire [15:0] reqs_1_bankEn = reqs_1_bankSel & _sourceD_wreq_out_bankEn_T_6; // @[BankedStore.scala 153:34]
  wire  regout_en = reqs_0_bankSel[0] | reqs_1_bankEn[0] | reqs_2_bankEn[0]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1 = reqs_1_bankSel[0]; // @[BankedStore.scala 180:33]
  wire  regout_wen = reqs_0_bankSel[0] | regout_sel_1; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T = regout_sel_1 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T = regout_sel_1 ? sourceD_wreq_words_0 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_0_io_r_req_valid_T = ~regout_wen; // @[BankedStore.scala 191:25]
  reg  regout_REG; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r; // @[Reg.scala 16:16]
  wire  regout_en_1 = reqs_0_bankSel[1] | reqs_1_bankEn[1] | reqs_2_bankEn[1]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_1 = reqs_1_bankSel[1]; // @[BankedStore.scala 180:33]
  wire  regout_wen_1 = reqs_0_bankSel[1] | regout_sel_1_1; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_1 = regout_sel_1_1 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_1 = regout_sel_1_1 ? sourceD_wreq_words_1 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_1_io_r_req_valid_T = ~regout_wen_1; // @[BankedStore.scala 191:25]
  reg  regout_REG_1; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_1; // @[Reg.scala 16:16]
  wire  regout_en_2 = reqs_0_bankSel[2] | reqs_1_bankEn[2] | reqs_2_bankEn[2]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_2 = reqs_1_bankSel[2]; // @[BankedStore.scala 180:33]
  wire  regout_wen_2 = reqs_0_bankSel[2] | regout_sel_1_2; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_2 = regout_sel_1_2 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_2 = regout_sel_1_2 ? sourceD_wreq_words_2 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_2_io_r_req_valid_T = ~regout_wen_2; // @[BankedStore.scala 191:25]
  reg  regout_REG_2; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_2; // @[Reg.scala 16:16]
  wire  regout_en_3 = reqs_0_bankSel[3] | reqs_1_bankEn[3] | reqs_2_bankEn[3]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_3 = reqs_1_bankSel[3]; // @[BankedStore.scala 180:33]
  wire  regout_wen_3 = reqs_0_bankSel[3] | regout_sel_1_3; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_3 = regout_sel_1_3 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_3 = regout_sel_1_3 ? sourceD_wreq_words_3 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_3_io_r_req_valid_T = ~regout_wen_3; // @[BankedStore.scala 191:25]
  reg  regout_REG_3; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_3; // @[Reg.scala 16:16]
  wire  regout_en_4 = reqs_0_bankSel[4] | reqs_1_bankEn[4] | reqs_2_bankEn[4]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_4 = reqs_1_bankSel[4]; // @[BankedStore.scala 180:33]
  wire  regout_wen_4 = reqs_0_bankSel[4] | regout_sel_1_4; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_4 = regout_sel_1_4 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_4 = regout_sel_1_4 ? sourceD_wreq_words_4 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_4_io_r_req_valid_T = ~regout_wen_4; // @[BankedStore.scala 191:25]
  reg  regout_REG_4; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_4; // @[Reg.scala 16:16]
  wire  regout_en_5 = reqs_0_bankSel[5] | reqs_1_bankEn[5] | reqs_2_bankEn[5]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_5 = reqs_1_bankSel[5]; // @[BankedStore.scala 180:33]
  wire  regout_wen_5 = reqs_0_bankSel[5] | regout_sel_1_5; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_5 = regout_sel_1_5 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_5 = regout_sel_1_5 ? sourceD_wreq_words_5 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_5_io_r_req_valid_T = ~regout_wen_5; // @[BankedStore.scala 191:25]
  reg  regout_REG_5; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_5; // @[Reg.scala 16:16]
  wire  regout_en_6 = reqs_0_bankSel[6] | reqs_1_bankEn[6] | reqs_2_bankEn[6]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_6 = reqs_1_bankSel[6]; // @[BankedStore.scala 180:33]
  wire  regout_wen_6 = reqs_0_bankSel[6] | regout_sel_1_6; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_6 = regout_sel_1_6 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_6 = regout_sel_1_6 ? sourceD_wreq_words_6 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_6_io_r_req_valid_T = ~regout_wen_6; // @[BankedStore.scala 191:25]
  reg  regout_REG_6; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_6; // @[Reg.scala 16:16]
  wire  regout_en_7 = reqs_0_bankSel[7] | reqs_1_bankEn[7] | reqs_2_bankEn[7]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_7 = reqs_1_bankSel[7]; // @[BankedStore.scala 180:33]
  wire  regout_wen_7 = reqs_0_bankSel[7] | regout_sel_1_7; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_7 = regout_sel_1_7 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_7 = regout_sel_1_7 ? sourceD_wreq_words_7 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_7_io_r_req_valid_T = ~regout_wen_7; // @[BankedStore.scala 191:25]
  reg  regout_REG_7; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_7; // @[Reg.scala 16:16]
  wire  regout_en_8 = reqs_0_bankSel[8] | reqs_1_bankEn[8] | reqs_2_bankEn[8]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_8 = reqs_1_bankSel[8]; // @[BankedStore.scala 180:33]
  wire  regout_wen_8 = reqs_0_bankSel[8] | regout_sel_1_8; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_8 = regout_sel_1_8 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_8 = regout_sel_1_8 ? sourceD_wreq_words_0 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_8_io_r_req_valid_T = ~regout_wen_8; // @[BankedStore.scala 191:25]
  reg  regout_REG_8; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_8; // @[Reg.scala 16:16]
  wire  regout_en_9 = reqs_0_bankSel[9] | reqs_1_bankEn[9] | reqs_2_bankEn[9]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_9 = reqs_1_bankSel[9]; // @[BankedStore.scala 180:33]
  wire  regout_wen_9 = reqs_0_bankSel[9] | regout_sel_1_9; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_9 = regout_sel_1_9 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_9 = regout_sel_1_9 ? sourceD_wreq_words_1 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_9_io_r_req_valid_T = ~regout_wen_9; // @[BankedStore.scala 191:25]
  reg  regout_REG_9; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_9; // @[Reg.scala 16:16]
  wire  regout_en_10 = reqs_0_bankSel[10] | reqs_1_bankEn[10] | reqs_2_bankEn[10]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_10 = reqs_1_bankSel[10]; // @[BankedStore.scala 180:33]
  wire  regout_wen_10 = reqs_0_bankSel[10] | regout_sel_1_10; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_10 = regout_sel_1_10 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_10 = regout_sel_1_10 ? sourceD_wreq_words_2 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_10_io_r_req_valid_T = ~regout_wen_10; // @[BankedStore.scala 191:25]
  reg  regout_REG_10; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_10; // @[Reg.scala 16:16]
  wire  regout_en_11 = reqs_0_bankSel[11] | reqs_1_bankEn[11] | reqs_2_bankEn[11]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_11 = reqs_1_bankSel[11]; // @[BankedStore.scala 180:33]
  wire  regout_wen_11 = reqs_0_bankSel[11] | regout_sel_1_11; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_11 = regout_sel_1_11 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_11 = regout_sel_1_11 ? sourceD_wreq_words_3 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_11_io_r_req_valid_T = ~regout_wen_11; // @[BankedStore.scala 191:25]
  reg  regout_REG_11; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_11; // @[Reg.scala 16:16]
  wire  regout_en_12 = reqs_0_bankSel[12] | reqs_1_bankEn[12] | reqs_2_bankEn[12]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_12 = reqs_1_bankSel[12]; // @[BankedStore.scala 180:33]
  wire  regout_wen_12 = reqs_0_bankSel[12] | regout_sel_1_12; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_12 = regout_sel_1_12 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_12 = regout_sel_1_12 ? sourceD_wreq_words_4 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_12_io_r_req_valid_T = ~regout_wen_12; // @[BankedStore.scala 191:25]
  reg  regout_REG_12; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_12; // @[Reg.scala 16:16]
  wire  regout_en_13 = reqs_0_bankSel[13] | reqs_1_bankEn[13] | reqs_2_bankEn[13]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_13 = reqs_1_bankSel[13]; // @[BankedStore.scala 180:33]
  wire  regout_wen_13 = reqs_0_bankSel[13] | regout_sel_1_13; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_13 = regout_sel_1_13 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_13 = regout_sel_1_13 ? sourceD_wreq_words_5 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_13_io_r_req_valid_T = ~regout_wen_13; // @[BankedStore.scala 191:25]
  reg  regout_REG_13; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_13; // @[Reg.scala 16:16]
  wire  regout_en_14 = reqs_0_bankSel[14] | reqs_1_bankEn[14] | reqs_2_bankEn[14]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_14 = reqs_1_bankSel[14]; // @[BankedStore.scala 180:33]
  wire  regout_wen_14 = reqs_0_bankSel[14] | regout_sel_1_14; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_14 = regout_sel_1_14 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_14 = regout_sel_1_14 ? sourceD_wreq_words_6 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_14_io_r_req_valid_T = ~regout_wen_14; // @[BankedStore.scala 191:25]
  reg  regout_REG_14; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_14; // @[Reg.scala 16:16]
  wire  regout_en_15 = reqs_0_bankSel[15] | reqs_1_bankEn[15] | reqs_2_bankEn[15]; // @[BankedStore.scala 179:45]
  wire  regout_sel_1_15 = reqs_1_bankSel[15]; // @[BankedStore.scala 180:33]
  wire  regout_wen_15 = reqs_0_bankSel[15] | regout_sel_1_15; // @[Mux.scala 47:70]
  wire [1:0] _regout_idx_T_15 = regout_sel_1_15 ? reqs_1_index : reqs_2_index; // @[Mux.scala 47:70]
  wire [31:0] _regout_data_T_15 = regout_sel_1_15 ? sourceD_wreq_words_7 : 32'h0; // @[Mux.scala 47:70]
  wire  _regout_cc_banks_15_io_r_req_valid_T = ~regout_wen_15; // @[BankedStore.scala 191:25]
  reg  regout_REG_15; // @[BankedStore.scala 193:43]
  reg [31:0] regout_r_15; // @[Reg.scala 16:16]
  reg [15:0] regsel_sourceD_REG; // @[BankedStore.scala 196:39]
  reg [15:0] regsel_sourceD; // @[BankedStore.scala 196:31]
  wire [31:0] _decodeDX_T_1 = regsel_sourceD[0] ? regout_r : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_3 = regsel_sourceD[1] ? regout_r_1 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_5 = regsel_sourceD[2] ? regout_r_2 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_7 = regsel_sourceD[3] ? regout_r_3 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_9 = regsel_sourceD[4] ? regout_r_4 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_11 = regsel_sourceD[5] ? regout_r_5 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_13 = regsel_sourceD[6] ? regout_r_6 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_15 = regsel_sourceD[7] ? regout_r_7 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_17 = regsel_sourceD[8] ? regout_r_8 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_19 = regsel_sourceD[9] ? regout_r_9 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_21 = regsel_sourceD[10] ? regout_r_10 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_23 = regsel_sourceD[11] ? regout_r_11 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_25 = regsel_sourceD[12] ? regout_r_12 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_27 = regsel_sourceD[13] ? regout_r_13 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_29 = regsel_sourceD[14] ? regout_r_14 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] _decodeDX_T_31 = regsel_sourceD[15] ? regout_r_15 : 32'h0; // @[BankedStore.scala 202:23]
  wire [31:0] decodeDX_0 = _decodeDX_T_1 | _decodeDX_T_17; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_1 = _decodeDX_T_3 | _decodeDX_T_19; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_2 = _decodeDX_T_5 | _decodeDX_T_21; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_3 = _decodeDX_T_7 | _decodeDX_T_23; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_4 = _decodeDX_T_9 | _decodeDX_T_25; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_5 = _decodeDX_T_11 | _decodeDX_T_27; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_6 = _decodeDX_T_13 | _decodeDX_T_29; // @[BankedStore.scala 203:85]
  wire [31:0] decodeDX_7 = _decodeDX_T_15 | _decodeDX_T_31; // @[BankedStore.scala 203:85]
  wire [127:0] io_sourceD_rdat_data_lo = {decodeDX_3,decodeDX_2,decodeDX_1,decodeDX_0}; // @[Cat.scala 31:58]
  wire [127:0] io_sourceD_rdat_data_hi = {decodeDX_7,decodeDX_6,decodeDX_5,decodeDX_4}; // @[Cat.scala 31:58]
  SRAMTemplate_39 cc_banks_0 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_0_clock),
    .reset(cc_banks_0_reset),
    .io_r_req_valid(cc_banks_0_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_0_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_0_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_0_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_0_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_0_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_1 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_1_clock),
    .reset(cc_banks_1_reset),
    .io_r_req_valid(cc_banks_1_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_1_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_1_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_1_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_1_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_1_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_2 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_2_clock),
    .reset(cc_banks_2_reset),
    .io_r_req_valid(cc_banks_2_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_2_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_2_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_2_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_2_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_2_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_3 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_3_clock),
    .reset(cc_banks_3_reset),
    .io_r_req_valid(cc_banks_3_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_3_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_3_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_3_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_3_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_3_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_4 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_4_clock),
    .reset(cc_banks_4_reset),
    .io_r_req_valid(cc_banks_4_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_4_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_4_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_4_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_4_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_4_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_5 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_5_clock),
    .reset(cc_banks_5_reset),
    .io_r_req_valid(cc_banks_5_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_5_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_5_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_5_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_5_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_5_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_6 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_6_clock),
    .reset(cc_banks_6_reset),
    .io_r_req_valid(cc_banks_6_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_6_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_6_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_6_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_6_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_6_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_7 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_7_clock),
    .reset(cc_banks_7_reset),
    .io_r_req_valid(cc_banks_7_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_7_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_7_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_7_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_7_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_7_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_8 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_8_clock),
    .reset(cc_banks_8_reset),
    .io_r_req_valid(cc_banks_8_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_8_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_8_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_8_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_8_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_8_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_9 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_9_clock),
    .reset(cc_banks_9_reset),
    .io_r_req_valid(cc_banks_9_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_9_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_9_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_9_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_9_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_9_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_10 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_10_clock),
    .reset(cc_banks_10_reset),
    .io_r_req_valid(cc_banks_10_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_10_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_10_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_10_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_10_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_10_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_11 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_11_clock),
    .reset(cc_banks_11_reset),
    .io_r_req_valid(cc_banks_11_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_11_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_11_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_11_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_11_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_11_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_12 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_12_clock),
    .reset(cc_banks_12_reset),
    .io_r_req_valid(cc_banks_12_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_12_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_12_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_12_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_12_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_12_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_13 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_13_clock),
    .reset(cc_banks_13_reset),
    .io_r_req_valid(cc_banks_13_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_13_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_13_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_13_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_13_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_13_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_14 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_14_clock),
    .reset(cc_banks_14_reset),
    .io_r_req_valid(cc_banks_14_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_14_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_14_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_14_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_14_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_14_io_w_req_bits_data_0)
  );
  SRAMTemplate_39 cc_banks_15 ( // @[BankedStore.scala 101:13]
    .clock(cc_banks_15_clock),
    .reset(cc_banks_15_reset),
    .io_r_req_valid(cc_banks_15_io_r_req_valid),
    .io_r_req_bits_setIdx(cc_banks_15_io_r_req_bits_setIdx),
    .io_r_resp_data_0(cc_banks_15_io_r_resp_data_0),
    .io_w_req_valid(cc_banks_15_io_w_req_valid),
    .io_w_req_bits_setIdx(cc_banks_15_io_w_req_bits_setIdx),
    .io_w_req_bits_data_0(cc_banks_15_io_w_req_bits_data_0)
  );
  assign io_sourceD_rdat_data = {io_sourceD_rdat_data_hi,io_sourceD_rdat_data_lo}; // @[Cat.scala 31:58]
  assign cc_banks_0_clock = clock;
  assign cc_banks_0_reset = reset;
  assign cc_banks_0_io_r_req_valid = ~regout_wen & regout_en; // @[BankedStore.scala 191:30]
  assign cc_banks_0_io_r_req_bits_setIdx = reqs_0_bankSel[0] ? reqs_0_index : _regout_idx_T; // @[Mux.scala 47:70]
  assign cc_banks_0_io_w_req_valid = regout_wen & regout_en; // @[BankedStore.scala 185:29]
  assign cc_banks_0_io_w_req_bits_setIdx = reqs_0_bankSel[0] ? reqs_0_index : _regout_idx_T; // @[Mux.scala 47:70]
  assign cc_banks_0_io_w_req_bits_data_0 = reqs_0_bankSel[0] ? sinkD_req_words_0 : _regout_data_T; // @[Mux.scala 47:70]
  assign cc_banks_1_clock = clock;
  assign cc_banks_1_reset = reset;
  assign cc_banks_1_io_r_req_valid = ~regout_wen_1 & regout_en_1; // @[BankedStore.scala 191:30]
  assign cc_banks_1_io_r_req_bits_setIdx = reqs_0_bankSel[1] ? reqs_0_index : _regout_idx_T_1; // @[Mux.scala 47:70]
  assign cc_banks_1_io_w_req_valid = regout_wen_1 & regout_en_1; // @[BankedStore.scala 185:29]
  assign cc_banks_1_io_w_req_bits_setIdx = reqs_0_bankSel[1] ? reqs_0_index : _regout_idx_T_1; // @[Mux.scala 47:70]
  assign cc_banks_1_io_w_req_bits_data_0 = reqs_0_bankSel[1] ? sinkD_req_words_1 : _regout_data_T_1; // @[Mux.scala 47:70]
  assign cc_banks_2_clock = clock;
  assign cc_banks_2_reset = reset;
  assign cc_banks_2_io_r_req_valid = ~regout_wen_2 & regout_en_2; // @[BankedStore.scala 191:30]
  assign cc_banks_2_io_r_req_bits_setIdx = reqs_0_bankSel[2] ? reqs_0_index : _regout_idx_T_2; // @[Mux.scala 47:70]
  assign cc_banks_2_io_w_req_valid = regout_wen_2 & regout_en_2; // @[BankedStore.scala 185:29]
  assign cc_banks_2_io_w_req_bits_setIdx = reqs_0_bankSel[2] ? reqs_0_index : _regout_idx_T_2; // @[Mux.scala 47:70]
  assign cc_banks_2_io_w_req_bits_data_0 = reqs_0_bankSel[2] ? sinkD_req_words_2 : _regout_data_T_2; // @[Mux.scala 47:70]
  assign cc_banks_3_clock = clock;
  assign cc_banks_3_reset = reset;
  assign cc_banks_3_io_r_req_valid = ~regout_wen_3 & regout_en_3; // @[BankedStore.scala 191:30]
  assign cc_banks_3_io_r_req_bits_setIdx = reqs_0_bankSel[3] ? reqs_0_index : _regout_idx_T_3; // @[Mux.scala 47:70]
  assign cc_banks_3_io_w_req_valid = regout_wen_3 & regout_en_3; // @[BankedStore.scala 185:29]
  assign cc_banks_3_io_w_req_bits_setIdx = reqs_0_bankSel[3] ? reqs_0_index : _regout_idx_T_3; // @[Mux.scala 47:70]
  assign cc_banks_3_io_w_req_bits_data_0 = reqs_0_bankSel[3] ? sinkD_req_words_3 : _regout_data_T_3; // @[Mux.scala 47:70]
  assign cc_banks_4_clock = clock;
  assign cc_banks_4_reset = reset;
  assign cc_banks_4_io_r_req_valid = ~regout_wen_4 & regout_en_4; // @[BankedStore.scala 191:30]
  assign cc_banks_4_io_r_req_bits_setIdx = reqs_0_bankSel[4] ? reqs_0_index : _regout_idx_T_4; // @[Mux.scala 47:70]
  assign cc_banks_4_io_w_req_valid = regout_wen_4 & regout_en_4; // @[BankedStore.scala 185:29]
  assign cc_banks_4_io_w_req_bits_setIdx = reqs_0_bankSel[4] ? reqs_0_index : _regout_idx_T_4; // @[Mux.scala 47:70]
  assign cc_banks_4_io_w_req_bits_data_0 = reqs_0_bankSel[4] ? sinkD_req_words_4 : _regout_data_T_4; // @[Mux.scala 47:70]
  assign cc_banks_5_clock = clock;
  assign cc_banks_5_reset = reset;
  assign cc_banks_5_io_r_req_valid = ~regout_wen_5 & regout_en_5; // @[BankedStore.scala 191:30]
  assign cc_banks_5_io_r_req_bits_setIdx = reqs_0_bankSel[5] ? reqs_0_index : _regout_idx_T_5; // @[Mux.scala 47:70]
  assign cc_banks_5_io_w_req_valid = regout_wen_5 & regout_en_5; // @[BankedStore.scala 185:29]
  assign cc_banks_5_io_w_req_bits_setIdx = reqs_0_bankSel[5] ? reqs_0_index : _regout_idx_T_5; // @[Mux.scala 47:70]
  assign cc_banks_5_io_w_req_bits_data_0 = reqs_0_bankSel[5] ? sinkD_req_words_5 : _regout_data_T_5; // @[Mux.scala 47:70]
  assign cc_banks_6_clock = clock;
  assign cc_banks_6_reset = reset;
  assign cc_banks_6_io_r_req_valid = ~regout_wen_6 & regout_en_6; // @[BankedStore.scala 191:30]
  assign cc_banks_6_io_r_req_bits_setIdx = reqs_0_bankSel[6] ? reqs_0_index : _regout_idx_T_6; // @[Mux.scala 47:70]
  assign cc_banks_6_io_w_req_valid = regout_wen_6 & regout_en_6; // @[BankedStore.scala 185:29]
  assign cc_banks_6_io_w_req_bits_setIdx = reqs_0_bankSel[6] ? reqs_0_index : _regout_idx_T_6; // @[Mux.scala 47:70]
  assign cc_banks_6_io_w_req_bits_data_0 = reqs_0_bankSel[6] ? sinkD_req_words_6 : _regout_data_T_6; // @[Mux.scala 47:70]
  assign cc_banks_7_clock = clock;
  assign cc_banks_7_reset = reset;
  assign cc_banks_7_io_r_req_valid = ~regout_wen_7 & regout_en_7; // @[BankedStore.scala 191:30]
  assign cc_banks_7_io_r_req_bits_setIdx = reqs_0_bankSel[7] ? reqs_0_index : _regout_idx_T_7; // @[Mux.scala 47:70]
  assign cc_banks_7_io_w_req_valid = regout_wen_7 & regout_en_7; // @[BankedStore.scala 185:29]
  assign cc_banks_7_io_w_req_bits_setIdx = reqs_0_bankSel[7] ? reqs_0_index : _regout_idx_T_7; // @[Mux.scala 47:70]
  assign cc_banks_7_io_w_req_bits_data_0 = reqs_0_bankSel[7] ? sinkD_req_words_7 : _regout_data_T_7; // @[Mux.scala 47:70]
  assign cc_banks_8_clock = clock;
  assign cc_banks_8_reset = reset;
  assign cc_banks_8_io_r_req_valid = ~regout_wen_8 & regout_en_8; // @[BankedStore.scala 191:30]
  assign cc_banks_8_io_r_req_bits_setIdx = reqs_0_bankSel[8] ? reqs_0_index : _regout_idx_T_8; // @[Mux.scala 47:70]
  assign cc_banks_8_io_w_req_valid = regout_wen_8 & regout_en_8; // @[BankedStore.scala 185:29]
  assign cc_banks_8_io_w_req_bits_setIdx = reqs_0_bankSel[8] ? reqs_0_index : _regout_idx_T_8; // @[Mux.scala 47:70]
  assign cc_banks_8_io_w_req_bits_data_0 = reqs_0_bankSel[8] ? sinkD_req_words_0 : _regout_data_T_8; // @[Mux.scala 47:70]
  assign cc_banks_9_clock = clock;
  assign cc_banks_9_reset = reset;
  assign cc_banks_9_io_r_req_valid = ~regout_wen_9 & regout_en_9; // @[BankedStore.scala 191:30]
  assign cc_banks_9_io_r_req_bits_setIdx = reqs_0_bankSel[9] ? reqs_0_index : _regout_idx_T_9; // @[Mux.scala 47:70]
  assign cc_banks_9_io_w_req_valid = regout_wen_9 & regout_en_9; // @[BankedStore.scala 185:29]
  assign cc_banks_9_io_w_req_bits_setIdx = reqs_0_bankSel[9] ? reqs_0_index : _regout_idx_T_9; // @[Mux.scala 47:70]
  assign cc_banks_9_io_w_req_bits_data_0 = reqs_0_bankSel[9] ? sinkD_req_words_1 : _regout_data_T_9; // @[Mux.scala 47:70]
  assign cc_banks_10_clock = clock;
  assign cc_banks_10_reset = reset;
  assign cc_banks_10_io_r_req_valid = ~regout_wen_10 & regout_en_10; // @[BankedStore.scala 191:30]
  assign cc_banks_10_io_r_req_bits_setIdx = reqs_0_bankSel[10] ? reqs_0_index : _regout_idx_T_10; // @[Mux.scala 47:70]
  assign cc_banks_10_io_w_req_valid = regout_wen_10 & regout_en_10; // @[BankedStore.scala 185:29]
  assign cc_banks_10_io_w_req_bits_setIdx = reqs_0_bankSel[10] ? reqs_0_index : _regout_idx_T_10; // @[Mux.scala 47:70]
  assign cc_banks_10_io_w_req_bits_data_0 = reqs_0_bankSel[10] ? sinkD_req_words_2 : _regout_data_T_10; // @[Mux.scala 47:70]
  assign cc_banks_11_clock = clock;
  assign cc_banks_11_reset = reset;
  assign cc_banks_11_io_r_req_valid = ~regout_wen_11 & regout_en_11; // @[BankedStore.scala 191:30]
  assign cc_banks_11_io_r_req_bits_setIdx = reqs_0_bankSel[11] ? reqs_0_index : _regout_idx_T_11; // @[Mux.scala 47:70]
  assign cc_banks_11_io_w_req_valid = regout_wen_11 & regout_en_11; // @[BankedStore.scala 185:29]
  assign cc_banks_11_io_w_req_bits_setIdx = reqs_0_bankSel[11] ? reqs_0_index : _regout_idx_T_11; // @[Mux.scala 47:70]
  assign cc_banks_11_io_w_req_bits_data_0 = reqs_0_bankSel[11] ? sinkD_req_words_3 : _regout_data_T_11; // @[Mux.scala 47:70]
  assign cc_banks_12_clock = clock;
  assign cc_banks_12_reset = reset;
  assign cc_banks_12_io_r_req_valid = ~regout_wen_12 & regout_en_12; // @[BankedStore.scala 191:30]
  assign cc_banks_12_io_r_req_bits_setIdx = reqs_0_bankSel[12] ? reqs_0_index : _regout_idx_T_12; // @[Mux.scala 47:70]
  assign cc_banks_12_io_w_req_valid = regout_wen_12 & regout_en_12; // @[BankedStore.scala 185:29]
  assign cc_banks_12_io_w_req_bits_setIdx = reqs_0_bankSel[12] ? reqs_0_index : _regout_idx_T_12; // @[Mux.scala 47:70]
  assign cc_banks_12_io_w_req_bits_data_0 = reqs_0_bankSel[12] ? sinkD_req_words_4 : _regout_data_T_12; // @[Mux.scala 47:70]
  assign cc_banks_13_clock = clock;
  assign cc_banks_13_reset = reset;
  assign cc_banks_13_io_r_req_valid = ~regout_wen_13 & regout_en_13; // @[BankedStore.scala 191:30]
  assign cc_banks_13_io_r_req_bits_setIdx = reqs_0_bankSel[13] ? reqs_0_index : _regout_idx_T_13; // @[Mux.scala 47:70]
  assign cc_banks_13_io_w_req_valid = regout_wen_13 & regout_en_13; // @[BankedStore.scala 185:29]
  assign cc_banks_13_io_w_req_bits_setIdx = reqs_0_bankSel[13] ? reqs_0_index : _regout_idx_T_13; // @[Mux.scala 47:70]
  assign cc_banks_13_io_w_req_bits_data_0 = reqs_0_bankSel[13] ? sinkD_req_words_5 : _regout_data_T_13; // @[Mux.scala 47:70]
  assign cc_banks_14_clock = clock;
  assign cc_banks_14_reset = reset;
  assign cc_banks_14_io_r_req_valid = ~regout_wen_14 & regout_en_14; // @[BankedStore.scala 191:30]
  assign cc_banks_14_io_r_req_bits_setIdx = reqs_0_bankSel[14] ? reqs_0_index : _regout_idx_T_14; // @[Mux.scala 47:70]
  assign cc_banks_14_io_w_req_valid = regout_wen_14 & regout_en_14; // @[BankedStore.scala 185:29]
  assign cc_banks_14_io_w_req_bits_setIdx = reqs_0_bankSel[14] ? reqs_0_index : _regout_idx_T_14; // @[Mux.scala 47:70]
  assign cc_banks_14_io_w_req_bits_data_0 = reqs_0_bankSel[14] ? sinkD_req_words_6 : _regout_data_T_14; // @[Mux.scala 47:70]
  assign cc_banks_15_clock = clock;
  assign cc_banks_15_reset = reset;
  assign cc_banks_15_io_r_req_valid = ~regout_wen_15 & regout_en_15; // @[BankedStore.scala 191:30]
  assign cc_banks_15_io_r_req_bits_setIdx = reqs_0_bankSel[15] ? reqs_0_index : _regout_idx_T_15; // @[Mux.scala 47:70]
  assign cc_banks_15_io_w_req_valid = regout_wen_15 & regout_en_15; // @[BankedStore.scala 185:29]
  assign cc_banks_15_io_w_req_bits_setIdx = reqs_0_bankSel[15] ? reqs_0_index : _regout_idx_T_15; // @[Mux.scala 47:70]
  assign cc_banks_15_io_w_req_bits_data_0 = reqs_0_bankSel[15] ? sinkD_req_words_7 : _regout_data_T_15; // @[Mux.scala 47:70]
  always @(posedge clock) begin
    regout_REG <= _regout_cc_banks_0_io_r_req_valid_T & regout_en; // @[BankedStore.scala 193:49]
    if (regout_REG) begin // @[Reg.scala 17:18]
      regout_r <= cc_banks_0_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_1 <= _regout_cc_banks_1_io_r_req_valid_T & regout_en_1; // @[BankedStore.scala 193:49]
    if (regout_REG_1) begin // @[Reg.scala 17:18]
      regout_r_1 <= cc_banks_1_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_2 <= _regout_cc_banks_2_io_r_req_valid_T & regout_en_2; // @[BankedStore.scala 193:49]
    if (regout_REG_2) begin // @[Reg.scala 17:18]
      regout_r_2 <= cc_banks_2_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_3 <= _regout_cc_banks_3_io_r_req_valid_T & regout_en_3; // @[BankedStore.scala 193:49]
    if (regout_REG_3) begin // @[Reg.scala 17:18]
      regout_r_3 <= cc_banks_3_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_4 <= _regout_cc_banks_4_io_r_req_valid_T & regout_en_4; // @[BankedStore.scala 193:49]
    if (regout_REG_4) begin // @[Reg.scala 17:18]
      regout_r_4 <= cc_banks_4_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_5 <= _regout_cc_banks_5_io_r_req_valid_T & regout_en_5; // @[BankedStore.scala 193:49]
    if (regout_REG_5) begin // @[Reg.scala 17:18]
      regout_r_5 <= cc_banks_5_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_6 <= _regout_cc_banks_6_io_r_req_valid_T & regout_en_6; // @[BankedStore.scala 193:49]
    if (regout_REG_6) begin // @[Reg.scala 17:18]
      regout_r_6 <= cc_banks_6_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_7 <= _regout_cc_banks_7_io_r_req_valid_T & regout_en_7; // @[BankedStore.scala 193:49]
    if (regout_REG_7) begin // @[Reg.scala 17:18]
      regout_r_7 <= cc_banks_7_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_8 <= _regout_cc_banks_8_io_r_req_valid_T & regout_en_8; // @[BankedStore.scala 193:49]
    if (regout_REG_8) begin // @[Reg.scala 17:18]
      regout_r_8 <= cc_banks_8_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_9 <= _regout_cc_banks_9_io_r_req_valid_T & regout_en_9; // @[BankedStore.scala 193:49]
    if (regout_REG_9) begin // @[Reg.scala 17:18]
      regout_r_9 <= cc_banks_9_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_10 <= _regout_cc_banks_10_io_r_req_valid_T & regout_en_10; // @[BankedStore.scala 193:49]
    if (regout_REG_10) begin // @[Reg.scala 17:18]
      regout_r_10 <= cc_banks_10_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_11 <= _regout_cc_banks_11_io_r_req_valid_T & regout_en_11; // @[BankedStore.scala 193:49]
    if (regout_REG_11) begin // @[Reg.scala 17:18]
      regout_r_11 <= cc_banks_11_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_12 <= _regout_cc_banks_12_io_r_req_valid_T & regout_en_12; // @[BankedStore.scala 193:49]
    if (regout_REG_12) begin // @[Reg.scala 17:18]
      regout_r_12 <= cc_banks_12_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_13 <= _regout_cc_banks_13_io_r_req_valid_T & regout_en_13; // @[BankedStore.scala 193:49]
    if (regout_REG_13) begin // @[Reg.scala 17:18]
      regout_r_13 <= cc_banks_13_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_14 <= _regout_cc_banks_14_io_r_req_valid_T & regout_en_14; // @[BankedStore.scala 193:49]
    if (regout_REG_14) begin // @[Reg.scala 17:18]
      regout_r_14 <= cc_banks_14_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regout_REG_15 <= _regout_cc_banks_15_io_r_req_valid_T & regout_en_15; // @[BankedStore.scala 193:49]
    if (regout_REG_15) begin // @[Reg.scala 17:18]
      regout_r_15 <= cc_banks_15_io_r_resp_data_0; // @[Reg.scala 17:22]
    end
    regsel_sourceD_REG <= reqs_2_bankSel & _sourceD_rreq_out_bankEn_T_6; // @[BankedStore.scala 153:34]
    regsel_sourceD <= regsel_sourceD_REG; // @[BankedStore.scala 196:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regout_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  regout_r = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regout_REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  regout_r_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regout_REG_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regout_r_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regout_REG_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  regout_r_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regout_REG_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  regout_r_4 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regout_REG_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  regout_r_5 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regout_REG_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  regout_r_6 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regout_REG_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  regout_r_7 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regout_REG_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  regout_r_8 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regout_REG_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  regout_r_9 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regout_REG_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  regout_r_10 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regout_REG_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  regout_r_11 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regout_REG_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  regout_r_12 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regout_REG_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  regout_r_13 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regout_REG_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  regout_r_14 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regout_REG_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  regout_r_15 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  regsel_sourceD_REG = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  regsel_sourceD = _RAND_33[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ListBuffer_1(
  input        clock,
  input        reset,
  output       io_push_ready,
  input        io_push_valid,
  input  [1:0] io_push_bits_index,
  input  [3:0] io_push_bits_data,
  output [3:0] io_valid,
  input        io_pop_valid,
  input  [1:0] io_pop_bits,
  output [3:0] io_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] head [0:3]; // @[ListBuffer.scala 51:18]
  wire  head_pop_head_en; // @[ListBuffer.scala 51:18]
  wire [1:0] head_pop_head_addr; // @[ListBuffer.scala 51:18]
  wire [1:0] head_pop_head_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_2_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_2_addr; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_2_mask; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_2_en; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_6_data; // @[ListBuffer.scala 51:18]
  wire [1:0] head_MPORT_6_addr; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_6_mask; // @[ListBuffer.scala 51:18]
  wire  head_MPORT_6_en; // @[ListBuffer.scala 51:18]
  reg [1:0] tail [0:3]; // @[ListBuffer.scala 52:18]
  wire  tail_push_tail_en; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_push_tail_addr; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_push_tail_data; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_4_en; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_4_addr; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_4_data; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_3_data; // @[ListBuffer.scala 52:18]
  wire [1:0] tail_MPORT_3_addr; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_3_mask; // @[ListBuffer.scala 52:18]
  wire  tail_MPORT_3_en; // @[ListBuffer.scala 52:18]
  reg [1:0] next [0:3]; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_5_en; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_5_addr; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_5_data; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_1_data; // @[ListBuffer.scala 54:18]
  wire [1:0] next_MPORT_1_addr; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_1_mask; // @[ListBuffer.scala 54:18]
  wire  next_MPORT_1_en; // @[ListBuffer.scala 54:18]
  reg [3:0] data [0:3]; // @[ListBuffer.scala 55:18]
  wire  data_io_data_MPORT_en; // @[ListBuffer.scala 55:18]
  wire [1:0] data_io_data_MPORT_addr; // @[ListBuffer.scala 55:18]
  wire [3:0] data_io_data_MPORT_data; // @[ListBuffer.scala 55:18]
  wire [3:0] data_MPORT_data; // @[ListBuffer.scala 55:18]
  wire [1:0] data_MPORT_addr; // @[ListBuffer.scala 55:18]
  wire  data_MPORT_mask; // @[ListBuffer.scala 55:18]
  wire  data_MPORT_en; // @[ListBuffer.scala 55:18]
  reg [3:0] valid; // @[ListBuffer.scala 50:22]
  reg [3:0] used; // @[ListBuffer.scala 53:22]
  wire [3:0] _freeOH_T = ~used; // @[ListBuffer.scala 57:27]
  wire [4:0] _freeOH_T_1 = {_freeOH_T, 1'h0}; // @[package.scala 244:48]
  wire [3:0] _freeOH_T_3 = _freeOH_T | _freeOH_T_1[3:0]; // @[package.scala 244:43]
  wire [5:0] _freeOH_T_4 = {_freeOH_T_3, 2'h0}; // @[package.scala 244:48]
  wire [3:0] _freeOH_T_6 = _freeOH_T_3 | _freeOH_T_4[3:0]; // @[package.scala 244:43]
  wire [4:0] _freeOH_T_8 = {_freeOH_T_6, 1'h0}; // @[ListBuffer.scala 57:44]
  wire [4:0] _freeOH_T_9 = ~_freeOH_T_8; // @[ListBuffer.scala 57:17]
  wire [4:0] _GEN_40 = {{1'd0}, _freeOH_T}; // @[ListBuffer.scala 57:60]
  wire [4:0] freeOH = _freeOH_T_9 & _GEN_40; // @[ListBuffer.scala 57:60]
  wire  freeIdx_hi = freeOH[4]; // @[OneHot.scala 30:18]
  wire [3:0] freeIdx_lo = freeOH[3:0]; // @[OneHot.scala 31:18]
  wire  _freeIdx_T = |freeIdx_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_41 = {{3'd0}, freeIdx_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _freeIdx_T_1 = _GEN_41 | freeIdx_lo; // @[OneHot.scala 32:28]
  wire [1:0] freeIdx_hi_1 = _freeIdx_T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] freeIdx_lo_1 = _freeIdx_T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _freeIdx_T_2 = |freeIdx_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _freeIdx_T_3 = freeIdx_hi_1 | freeIdx_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] freeIdx = {_freeIdx_T,_freeIdx_T_2,_freeIdx_T_3[1]}; // @[Cat.scala 31:58]
  wire [3:0] _push_valid_T = valid >> io_push_bits_index; // @[ListBuffer.scala 70:25]
  wire  push_valid = _push_valid_T[0]; // @[ListBuffer.scala 70:25]
  wire  _T = io_push_ready & io_push_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _valid_set_T = 4'h1 << io_push_bits_index; // @[OneHot.scala 64:12]
  wire  _GEN_7 = push_valid ? 1'h0 : 1'h1; // @[ListBuffer.scala 51:18 77:23]
  wire [3:0] valid_set = _T ? _valid_set_T : 4'h0; // @[ListBuffer.scala 73:25 74:15]
  wire [4:0] _GEN_11 = _T ? freeOH : 5'h0; // @[ListBuffer.scala 73:25 75:14]
  wire  _GEN_19 = _T & push_valid; // @[ListBuffer.scala 54:18 73:25]
  wire [3:0] _T_3 = io_valid >> io_pop_bits; // @[ListBuffer.scala 101:39]
  wire [1:0] used_clr_shiftAmount = head_pop_head_data; // @[OneHot.scala 63:49]
  wire [3:0] _used_clr_T = 4'h1 << used_clr_shiftAmount; // @[OneHot.scala 64:12]
  wire [3:0] _valid_clr_T = 4'h1 << io_pop_bits; // @[OneHot.scala 64:12]
  wire [3:0] _GEN_29 = head_pop_head_data == tail_MPORT_4_data ? _valid_clr_T : 4'h0; // @[ListBuffer.scala 108:48 109:17]
  wire [2:0] _T_14 = _GEN_19 & tail_push_tail_data == head_pop_head_data ? freeIdx : {{1'd0}, next_MPORT_5_data}; // @[ListBuffer.scala 111:32]
  wire [3:0] used_clr = io_pop_valid ? _used_clr_T : 4'h0; // @[ListBuffer.scala 106:24 107:14]
  wire [3:0] valid_clr = io_pop_valid ? _GEN_29 : 4'h0; // @[ListBuffer.scala 106:24]
  wire [3:0] _used_T = ~used_clr; // @[ListBuffer.scala 124:24]
  wire [3:0] _used_T_1 = used & _used_T; // @[ListBuffer.scala 124:21]
  wire [3:0] used_set = _GEN_11[3:0];
  wire [3:0] _used_T_4 = _used_T_1 | used_set; // @[ListBuffer.scala 124:70]
  wire [3:0] _valid_T = ~valid_clr; // @[ListBuffer.scala 125:24]
  wire [3:0] _valid_T_1 = valid & _valid_T; // @[ListBuffer.scala 125:21]
  wire [3:0] _valid_T_4 = _valid_T_1 | valid_set; // @[ListBuffer.scala 125:71]
  assign head_pop_head_en = 1'h1;
  assign head_pop_head_addr = io_pop_bits;
  assign head_pop_head_data = head[head_pop_head_addr]; // @[ListBuffer.scala 51:18]
  assign head_MPORT_2_data = freeIdx[1:0];
  assign head_MPORT_2_addr = io_push_bits_index;
  assign head_MPORT_2_mask = 1'h1;
  assign head_MPORT_2_en = _T & _GEN_7;
  assign head_MPORT_6_data = _T_14[1:0];
  assign head_MPORT_6_addr = io_pop_bits;
  assign head_MPORT_6_mask = 1'h1;
  assign head_MPORT_6_en = io_pop_valid;
  assign tail_push_tail_en = 1'h1;
  assign tail_push_tail_addr = io_push_bits_index;
  assign tail_push_tail_data = tail[tail_push_tail_addr]; // @[ListBuffer.scala 52:18]
  assign tail_MPORT_4_en = io_pop_valid;
  assign tail_MPORT_4_addr = io_pop_bits;
  assign tail_MPORT_4_data = tail[tail_MPORT_4_addr]; // @[ListBuffer.scala 52:18]
  assign tail_MPORT_3_data = freeIdx[1:0];
  assign tail_MPORT_3_addr = io_push_bits_index;
  assign tail_MPORT_3_mask = 1'h1;
  assign tail_MPORT_3_en = io_push_ready & io_push_valid;
  assign next_MPORT_5_en = io_pop_valid;
  assign next_MPORT_5_addr = head_pop_head_data;
  assign next_MPORT_5_data = next[next_MPORT_5_addr]; // @[ListBuffer.scala 54:18]
  assign next_MPORT_1_data = freeIdx[1:0];
  assign next_MPORT_1_addr = tail_push_tail_data;
  assign next_MPORT_1_mask = 1'h1;
  assign next_MPORT_1_en = _T & push_valid;
  assign data_io_data_MPORT_en = 1'h1;
  assign data_io_data_MPORT_addr = head_pop_head_data;
  assign data_io_data_MPORT_data = data[data_io_data_MPORT_addr]; // @[ListBuffer.scala 55:18]
  assign data_MPORT_data = io_push_bits_data;
  assign data_MPORT_addr = freeIdx[1:0];
  assign data_MPORT_mask = 1'h1;
  assign data_MPORT_en = io_push_ready & io_push_valid;
  assign io_push_ready = ~(&used); // @[ListBuffer.scala 72:20]
  assign io_valid = valid; // @[ListBuffer.scala 98:12]
  assign io_data = data_io_data_MPORT_data; // @[ListBuffer.scala 96:{63,63}]
  always @(posedge clock) begin
    if (head_MPORT_2_en & head_MPORT_2_mask) begin
      head[head_MPORT_2_addr] <= head_MPORT_2_data; // @[ListBuffer.scala 51:18]
    end
    if (head_MPORT_6_en & head_MPORT_6_mask) begin
      head[head_MPORT_6_addr] <= head_MPORT_6_data; // @[ListBuffer.scala 51:18]
    end
    if (tail_MPORT_3_en & tail_MPORT_3_mask) begin
      tail[tail_MPORT_3_addr] <= tail_MPORT_3_data; // @[ListBuffer.scala 52:18]
    end
    if (next_MPORT_1_en & next_MPORT_1_mask) begin
      next[next_MPORT_1_addr] <= next_MPORT_1_data; // @[ListBuffer.scala 54:18]
    end
    if (data_MPORT_en & data_MPORT_mask) begin
      data[data_MPORT_addr] <= data_MPORT_data; // @[ListBuffer.scala 55:18]
    end
    if (reset) begin // @[ListBuffer.scala 50:22]
      valid <= 4'h0; // @[ListBuffer.scala 50:22]
    end else begin
      valid <= _valid_T_4;
    end
    if (reset) begin // @[ListBuffer.scala 53:22]
      used <= 4'h0; // @[ListBuffer.scala 53:22]
    end else begin
      used <= _used_T_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(~io_pop_valid | _T_3[0])) begin
          $fatal; // @[ListBuffer.scala 101:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_pop_valid | _T_3[0])) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ListBuffer.scala:101 assert (!io.pop.fire() || (io.valid)(io.pop.bits))\n"); // @[ListBuffer.scala 101:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    head[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    tail[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    next[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    data[initvar] = _RAND_3[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  valid = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  used = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MSHR_4(
  input          clock,
  input          reset,
  input          io_allocate_valid,
  input  [2:0]   io_allocate_bits_opcode,
  input  [25:0]  io_allocate_bits_tag,
  input  [4:0]   io_allocate_bits_offset,
  input  [1:0]   io_allocate_bits_put,
  input  [255:0] io_allocate_bits_data,
  input  [7:0]   io_allocate_bits_mask,
  input          io_allocate_bits_set,
  input  [1:0]   io_allocate_bits_way,
  output [2:0]   io_status_opcode,
  output [25:0]  io_status_tag,
  output [1:0]   io_status_put,
  output         io_status_set,
  output [1:0]   io_status_way,
  input          io_valid,
  input          io_schedule_a_ready,
  output         io_schedule_a_valid,
  output [25:0]  io_schedule_a_bits_tag,
  output [4:0]   io_schedule_a_bits_offset,
  output [255:0] io_schedule_a_bits_data,
  output         io_schedule_a_bits_set,
  output         io_schedule_d_valid,
  output [2:0]   io_schedule_d_bits_opcode,
  output [25:0]  io_schedule_d_bits_tag,
  output [4:0]   io_schedule_d_bits_offset,
  output [1:0]   io_schedule_d_bits_put,
  output [255:0] io_schedule_d_bits_data,
  output [7:0]   io_schedule_d_bits_mask,
  output         io_schedule_d_bits_set,
  output [1:0]   io_schedule_d_bits_way,
  input          io_schedule_dir_ready,
  output         io_schedule_dir_valid,
  output [1:0]   io_schedule_dir_bits_way,
  output [25:0]  io_schedule_dir_bits_data_tag,
  output         io_schedule_dir_bits_set,
  input          io_sinkd_valid,
  input  [255:0] io_sinkd_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] request_opcode; // @[MSHR.scala 51:24]
  reg [25:0] request_tag; // @[MSHR.scala 51:24]
  reg [4:0] request_offset; // @[MSHR.scala 51:24]
  reg [1:0] request_put; // @[MSHR.scala 51:24]
  reg [255:0] request_data; // @[MSHR.scala 51:24]
  reg [7:0] request_mask; // @[MSHR.scala 51:24]
  reg  request_set; // @[MSHR.scala 51:24]
  reg [1:0] request_way; // @[MSHR.scala 51:24]
  reg  sche_a_valid; // @[MSHR.scala 62:27]
  reg  sche_dir_valid; // @[MSHR.scala 63:29]
  reg  sink_d_reg; // @[MSHR.scala 64:25]
  wire  _GEN_11 = io_allocate_valid ? 1'h0 : sink_d_reg; // @[MSHR.scala 66:28 68:15 64:25]
  wire  _T = io_schedule_a_ready & io_schedule_a_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = io_schedule_dir_ready & io_schedule_dir_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_13 = _T_1 ? 1'h0 : sche_dir_valid; // @[MSHR.scala 63:29 91:{31,46}]
  wire  _GEN_14 = io_sinkd_valid | _GEN_13; // @[MSHR.scala 104:25 105:19]
  wire  _GEN_15 = io_sinkd_valid | _GEN_11; // @[MSHR.scala 104:25 106:16]
  assign io_status_opcode = request_opcode; // @[MSHR.scala 57:16]
  assign io_status_tag = request_tag; // @[MSHR.scala 57:16]
  assign io_status_put = request_put; // @[MSHR.scala 57:16]
  assign io_status_set = request_set; // @[MSHR.scala 57:16]
  assign io_status_way = request_way; // @[MSHR.scala 57:16]
  assign io_schedule_a_valid = sche_a_valid; // @[MSHR.scala 79:22]
  assign io_schedule_a_bits_tag = request_tag; // @[MSHR.scala 82:25]
  assign io_schedule_a_bits_offset = request_offset; // @[MSHR.scala 84:28]
  assign io_schedule_a_bits_data = request_data; // @[MSHR.scala 86:26]
  assign io_schedule_a_bits_set = request_set; // @[MSHR.scala 80:25]
  assign io_schedule_d_valid = io_valid & sink_d_reg; // @[MSHR.scala 72:34]
  assign io_schedule_d_bits_opcode = request_opcode; // @[MSHR.scala 73:21]
  assign io_schedule_d_bits_tag = request_tag; // @[MSHR.scala 73:21]
  assign io_schedule_d_bits_offset = request_offset; // @[MSHR.scala 73:21]
  assign io_schedule_d_bits_put = request_put; // @[MSHR.scala 73:21]
  assign io_schedule_d_bits_data = sink_d_reg ? io_sinkd_bits_data : request_data; // @[MSHR.scala 75:32]
  assign io_schedule_d_bits_mask = request_mask; // @[MSHR.scala 73:21]
  assign io_schedule_d_bits_set = request_set; // @[MSHR.scala 73:21]
  assign io_schedule_d_bits_way = request_way; // @[MSHR.scala 73:21]
  assign io_schedule_dir_valid = sche_dir_valid; // @[MSHR.scala 94:24]
  assign io_schedule_dir_bits_way = request_way; // @[MSHR.scala 98:27]
  assign io_schedule_dir_bits_data_tag = request_tag; // @[MSHR.scala 96:32]
  assign io_schedule_dir_bits_set = request_set; // @[MSHR.scala 95:27]
  always @(posedge clock) begin
    if (reset) begin // @[MSHR.scala 51:24]
      request_opcode <= 3'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_opcode <= io_allocate_bits_opcode; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_tag <= 26'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_tag <= io_allocate_bits_tag; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_offset <= 5'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_offset <= io_allocate_bits_offset; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_put <= 2'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_put <= io_allocate_bits_put; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_data <= 256'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_data <= io_allocate_bits_data; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_mask <= 8'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_mask <= io_allocate_bits_mask; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_set <= 1'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_set <= io_allocate_bits_set; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 51:24]
      request_way <= 2'h0; // @[MSHR.scala 51:24]
    end else if (io_allocate_valid) begin // @[MSHR.scala 66:28]
      request_way <= io_allocate_bits_way; // @[MSHR.scala 67:13]
    end
    if (reset) begin // @[MSHR.scala 62:27]
      sche_a_valid <= 1'h0; // @[MSHR.scala 62:27]
    end else if (_T) begin // @[MSHR.scala 89:29]
      sche_a_valid <= 1'h0; // @[MSHR.scala 89:42]
    end else begin
      sche_a_valid <= io_allocate_valid; // @[MSHR.scala 78:15]
    end
    if (reset) begin // @[MSHR.scala 63:29]
      sche_dir_valid <= 1'h0; // @[MSHR.scala 63:29]
    end else begin
      sche_dir_valid <= _GEN_14;
    end
    if (reset) begin // @[MSHR.scala 64:25]
      sink_d_reg <= 1'h0; // @[MSHR.scala 64:25]
    end else begin
      sink_d_reg <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  request_opcode = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  request_tag = _RAND_1[25:0];
  _RAND_2 = {1{`RANDOM}};
  request_offset = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  request_put = _RAND_3[1:0];
  _RAND_4 = {8{`RANDOM}};
  request_data = _RAND_4[255:0];
  _RAND_5 = {1{`RANDOM}};
  request_mask = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  request_set = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  request_way = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  sche_a_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sche_dir_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sink_d_reg = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_106(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [3:0]   io_enq_bits_source,
  input  [25:0]  io_enq_bits_tag,
  input  [4:0]   io_enq_bits_offset,
  input  [255:0] io_enq_bits_data,
  input  [7:0]   io_enq_bits_mask,
  input          io_enq_bits_set,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [3:0]   io_deq_bits_source,
  output [25:0]  io_deq_bits_tag,
  output [4:0]   io_deq_bits_offset,
  output [255:0] io_deq_bits_data,
  output [7:0]   io_deq_bits_mask,
  output         io_deq_bits_set
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_source [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [25:0] ram_tag [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_tag_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [25:0] ram_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [25:0] ram_tag_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_tag_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_offset [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_offset_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_offset_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_offset_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_offset_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_offset_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_offset_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_offset_MPORT_en; // @[Decoupled.scala 259:95]
  reg [255:0] ram_data [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [255:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [255:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_set [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_set_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_set_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_set_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_set_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_set_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_set_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_set_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = 3'h0;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tag_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tag_io_deq_bits_MPORT_data = ram_tag[ram_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_tag_MPORT_data = io_enq_bits_tag;
  assign ram_tag_MPORT_addr = enq_ptr_value;
  assign ram_tag_MPORT_mask = 1'h1;
  assign ram_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_offset_io_deq_bits_MPORT_en = 1'h1;
  assign ram_offset_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_offset_io_deq_bits_MPORT_data = ram_offset[ram_offset_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_offset_MPORT_data = io_enq_bits_offset;
  assign ram_offset_MPORT_addr = enq_ptr_value;
  assign ram_offset_MPORT_mask = 1'h1;
  assign ram_offset_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_set_io_deq_bits_MPORT_en = 1'h1;
  assign ram_set_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_set_io_deq_bits_MPORT_data = ram_set[ram_set_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_set_MPORT_data = io_enq_bits_set;
  assign ram_set_MPORT_addr = enq_ptr_value;
  assign ram_set_MPORT_mask = 1'h1;
  assign ram_set_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_tag = ram_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_offset = ram_offset_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_set = ram_set_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_tag_MPORT_en & ram_tag_MPORT_mask) begin
      ram_tag[ram_tag_MPORT_addr] <= ram_tag_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_offset_MPORT_en & ram_offset_MPORT_mask) begin
      ram_offset[ram_offset_MPORT_addr] <= ram_offset_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_set_MPORT_en & ram_set_MPORT_mask) begin
      ram_set[ram_set_MPORT_addr] <= ram_set_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_source[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_tag[initvar] = _RAND_2[25:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_offset[initvar] = _RAND_3[4:0];
  _RAND_4 = {8{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[255:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_set[initvar] = _RAND_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enq_ptr_value = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  deq_ptr_value = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_107(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [2:0]   io_enq_bits_opcode,
  input  [3:0]   io_enq_bits_source,
  input  [25:0]  io_enq_bits_tag,
  input  [4:0]   io_enq_bits_offset,
  input  [1:0]   io_enq_bits_put,
  input  [255:0] io_enq_bits_data,
  input  [7:0]   io_enq_bits_mask,
  input          io_enq_bits_set,
  input          io_enq_bits_hit,
  input  [1:0]   io_enq_bits_way,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [3:0]   io_deq_bits_source,
  output [25:0]  io_deq_bits_tag,
  output [4:0]   io_deq_bits_offset,
  output [1:0]   io_deq_bits_put,
  output [255:0] io_deq_bits_data,
  output [7:0]   io_deq_bits_mask,
  output         io_deq_bits_set,
  output         io_deq_bits_hit,
  output [1:0]   io_deq_bits_way
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [255:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_source [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [25:0] ram_tag [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_tag_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [25:0] ram_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [25:0] ram_tag_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_tag_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_offset [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_offset_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_offset_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_offset_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_offset_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_offset_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_offset_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_offset_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_put [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_put_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_put_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_put_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_put_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_put_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_put_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_put_MPORT_en; // @[Decoupled.scala 259:95]
  reg [255:0] ram_data [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [255:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [255:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_set [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_set_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_set_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_set_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_set_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_set_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_set_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_set_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_hit [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_hit_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_hit_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_hit_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_hit_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_hit_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_hit_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_hit_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_way [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_way_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_way_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_way_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_way_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_way_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_way_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_way_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tag_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tag_io_deq_bits_MPORT_data = ram_tag[ram_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_tag_MPORT_data = io_enq_bits_tag;
  assign ram_tag_MPORT_addr = enq_ptr_value;
  assign ram_tag_MPORT_mask = 1'h1;
  assign ram_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_offset_io_deq_bits_MPORT_en = 1'h1;
  assign ram_offset_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_offset_io_deq_bits_MPORT_data = ram_offset[ram_offset_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_offset_MPORT_data = io_enq_bits_offset;
  assign ram_offset_MPORT_addr = enq_ptr_value;
  assign ram_offset_MPORT_mask = 1'h1;
  assign ram_offset_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_put_io_deq_bits_MPORT_en = 1'h1;
  assign ram_put_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_put_io_deq_bits_MPORT_data = ram_put[ram_put_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_put_MPORT_data = io_enq_bits_put;
  assign ram_put_MPORT_addr = enq_ptr_value;
  assign ram_put_MPORT_mask = 1'h1;
  assign ram_put_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_set_io_deq_bits_MPORT_en = 1'h1;
  assign ram_set_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_set_io_deq_bits_MPORT_data = ram_set[ram_set_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_set_MPORT_data = io_enq_bits_set;
  assign ram_set_MPORT_addr = enq_ptr_value;
  assign ram_set_MPORT_mask = 1'h1;
  assign ram_set_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_hit_io_deq_bits_MPORT_en = 1'h1;
  assign ram_hit_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_hit_io_deq_bits_MPORT_data = ram_hit[ram_hit_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_hit_MPORT_data = io_enq_bits_hit;
  assign ram_hit_MPORT_addr = enq_ptr_value;
  assign ram_hit_MPORT_mask = 1'h1;
  assign ram_hit_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_way_io_deq_bits_MPORT_en = 1'h1;
  assign ram_way_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_way_io_deq_bits_MPORT_data = ram_way[ram_way_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_way_MPORT_data = io_enq_bits_way;
  assign ram_way_MPORT_addr = enq_ptr_value;
  assign ram_way_MPORT_mask = 1'h1;
  assign ram_way_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_tag = ram_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_offset = ram_offset_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_put = ram_put_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_set = ram_set_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_hit = ram_hit_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_way = ram_way_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_tag_MPORT_en & ram_tag_MPORT_mask) begin
      ram_tag[ram_tag_MPORT_addr] <= ram_tag_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_offset_MPORT_en & ram_offset_MPORT_mask) begin
      ram_offset[ram_offset_MPORT_addr] <= ram_offset_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_put_MPORT_en & ram_put_MPORT_mask) begin
      ram_put[ram_put_MPORT_addr] <= ram_put_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_set_MPORT_en & ram_set_MPORT_mask) begin
      ram_set[ram_set_MPORT_addr] <= ram_set_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_hit_MPORT_en & ram_hit_MPORT_mask) begin
      ram_hit[ram_hit_MPORT_addr] <= ram_hit_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_way_MPORT_en & ram_way_MPORT_mask) begin
      ram_way[ram_way_MPORT_addr] <= ram_way_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_source[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_tag[initvar] = _RAND_2[25:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_offset[initvar] = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_put[initvar] = _RAND_4[1:0];
  _RAND_5 = {8{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[255:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_mask[initvar] = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_set[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_hit[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_way[initvar] = _RAND_9[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  enq_ptr_value = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  deq_ptr_value = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  maybe_full = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scheduler(
  input          clock,
  input          reset,
  output         io_in_a_ready,
  input          io_in_a_valid,
  input  [2:0]   io_in_a_bits_opcode,
  input  [3:0]   io_in_a_bits_source,
  input  [31:0]  io_in_a_bits_address,
  input  [31:0]  io_in_a_bits_mask,
  input  [255:0] io_in_a_bits_data,
  input          io_in_d_ready,
  output         io_in_d_valid,
  output [3:0]   io_in_d_bits_source,
  output [255:0] io_in_d_bits_data,
  output [31:0]  io_in_d_bits_address,
  input          io_out_a_ready,
  output         io_out_a_valid,
  output [2:0]   io_out_a_bits_opcode,
  output [3:0]   io_out_a_bits_source,
  output [31:0]  io_out_a_bits_address,
  output [31:0]  io_out_a_bits_mask,
  output [255:0] io_out_a_bits_data,
  output         io_out_d_ready,
  input          io_out_d_valid,
  input  [2:0]   io_out_d_bits_opcode,
  input  [3:0]   io_out_d_bits_source,
  input  [255:0] io_out_d_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  sourceA_io_req_ready; // @[Scheduler.scala 49:23]
  wire  sourceA_io_req_valid; // @[Scheduler.scala 49:23]
  wire [2:0] sourceA_io_req_bits_opcode; // @[Scheduler.scala 49:23]
  wire [3:0] sourceA_io_req_bits_source; // @[Scheduler.scala 49:23]
  wire [25:0] sourceA_io_req_bits_tag; // @[Scheduler.scala 49:23]
  wire [4:0] sourceA_io_req_bits_offset; // @[Scheduler.scala 49:23]
  wire [255:0] sourceA_io_req_bits_data; // @[Scheduler.scala 49:23]
  wire [7:0] sourceA_io_req_bits_mask; // @[Scheduler.scala 49:23]
  wire  sourceA_io_req_bits_set; // @[Scheduler.scala 49:23]
  wire  sourceA_io_a_ready; // @[Scheduler.scala 49:23]
  wire  sourceA_io_a_valid; // @[Scheduler.scala 49:23]
  wire [2:0] sourceA_io_a_bits_opcode; // @[Scheduler.scala 49:23]
  wire [3:0] sourceA_io_a_bits_source; // @[Scheduler.scala 49:23]
  wire [31:0] sourceA_io_a_bits_address; // @[Scheduler.scala 49:23]
  wire [31:0] sourceA_io_a_bits_mask; // @[Scheduler.scala 49:23]
  wire [255:0] sourceA_io_a_bits_data; // @[Scheduler.scala 49:23]
  wire  sourceD_clock; // @[Scheduler.scala 51:23]
  wire  sourceD_reset; // @[Scheduler.scala 51:23]
  wire  sourceD_io_req_ready; // @[Scheduler.scala 51:23]
  wire  sourceD_io_req_valid; // @[Scheduler.scala 51:23]
  wire [2:0] sourceD_io_req_bits_opcode; // @[Scheduler.scala 51:23]
  wire [3:0] sourceD_io_req_bits_source; // @[Scheduler.scala 51:23]
  wire [25:0] sourceD_io_req_bits_tag; // @[Scheduler.scala 51:23]
  wire [4:0] sourceD_io_req_bits_offset; // @[Scheduler.scala 51:23]
  wire [1:0] sourceD_io_req_bits_put; // @[Scheduler.scala 51:23]
  wire [255:0] sourceD_io_req_bits_data; // @[Scheduler.scala 51:23]
  wire [7:0] sourceD_io_req_bits_mask; // @[Scheduler.scala 51:23]
  wire  sourceD_io_req_bits_set; // @[Scheduler.scala 51:23]
  wire  sourceD_io_req_bits_hit; // @[Scheduler.scala 51:23]
  wire [1:0] sourceD_io_req_bits_way; // @[Scheduler.scala 51:23]
  wire  sourceD_io_req_bits_from_mem; // @[Scheduler.scala 51:23]
  wire  sourceD_io_d_ready; // @[Scheduler.scala 51:23]
  wire  sourceD_io_d_valid; // @[Scheduler.scala 51:23]
  wire [3:0] sourceD_io_d_bits_source; // @[Scheduler.scala 51:23]
  wire [255:0] sourceD_io_d_bits_data; // @[Scheduler.scala 51:23]
  wire [31:0] sourceD_io_d_bits_address; // @[Scheduler.scala 51:23]
  wire  sourceD_io_pb_pop_valid; // @[Scheduler.scala 51:23]
  wire [1:0] sourceD_io_pb_pop_bits_index; // @[Scheduler.scala 51:23]
  wire [255:0] sourceD_io_pb_beat_data; // @[Scheduler.scala 51:23]
  wire [7:0] sourceD_io_pb_beat_mask; // @[Scheduler.scala 51:23]
  wire  sourceD_io_bs_radr_valid; // @[Scheduler.scala 51:23]
  wire [1:0] sourceD_io_bs_radr_bits_way; // @[Scheduler.scala 51:23]
  wire  sourceD_io_bs_radr_bits_set; // @[Scheduler.scala 51:23]
  wire [7:0] sourceD_io_bs_radr_bits_mask; // @[Scheduler.scala 51:23]
  wire [255:0] sourceD_io_bs_rdat_data; // @[Scheduler.scala 51:23]
  wire  sourceD_io_bs_wadr_valid; // @[Scheduler.scala 51:23]
  wire [1:0] sourceD_io_bs_wadr_bits_way; // @[Scheduler.scala 51:23]
  wire  sourceD_io_bs_wadr_bits_set; // @[Scheduler.scala 51:23]
  wire [7:0] sourceD_io_bs_wadr_bits_mask; // @[Scheduler.scala 51:23]
  wire [255:0] sourceD_io_bs_wdat_data; // @[Scheduler.scala 51:23]
  wire  sourceD_io_a_ready; // @[Scheduler.scala 51:23]
  wire  sourceD_io_a_valid; // @[Scheduler.scala 51:23]
  wire [3:0] sourceD_io_a_bits_source; // @[Scheduler.scala 51:23]
  wire [25:0] sourceD_io_a_bits_tag; // @[Scheduler.scala 51:23]
  wire [4:0] sourceD_io_a_bits_offset; // @[Scheduler.scala 51:23]
  wire [255:0] sourceD_io_a_bits_data; // @[Scheduler.scala 51:23]
  wire [7:0] sourceD_io_a_bits_mask; // @[Scheduler.scala 51:23]
  wire  sourceD_io_a_bits_set; // @[Scheduler.scala 51:23]
  wire  sinkA_clock; // @[Scheduler.scala 53:21]
  wire  sinkA_reset; // @[Scheduler.scala 53:21]
  wire  sinkA_io_req_ready; // @[Scheduler.scala 53:21]
  wire  sinkA_io_req_valid; // @[Scheduler.scala 53:21]
  wire [2:0] sinkA_io_req_bits_opcode; // @[Scheduler.scala 53:21]
  wire [3:0] sinkA_io_req_bits_source; // @[Scheduler.scala 53:21]
  wire [25:0] sinkA_io_req_bits_tag; // @[Scheduler.scala 53:21]
  wire [4:0] sinkA_io_req_bits_offset; // @[Scheduler.scala 53:21]
  wire [1:0] sinkA_io_req_bits_put; // @[Scheduler.scala 53:21]
  wire [255:0] sinkA_io_req_bits_data; // @[Scheduler.scala 53:21]
  wire [7:0] sinkA_io_req_bits_mask; // @[Scheduler.scala 53:21]
  wire  sinkA_io_req_bits_set; // @[Scheduler.scala 53:21]
  wire  sinkA_io_a_ready; // @[Scheduler.scala 53:21]
  wire  sinkA_io_a_valid; // @[Scheduler.scala 53:21]
  wire [2:0] sinkA_io_a_bits_opcode; // @[Scheduler.scala 53:21]
  wire [3:0] sinkA_io_a_bits_source; // @[Scheduler.scala 53:21]
  wire [31:0] sinkA_io_a_bits_address; // @[Scheduler.scala 53:21]
  wire [31:0] sinkA_io_a_bits_mask; // @[Scheduler.scala 53:21]
  wire [255:0] sinkA_io_a_bits_data; // @[Scheduler.scala 53:21]
  wire  sinkA_io_pb_pop_ready; // @[Scheduler.scala 53:21]
  wire  sinkA_io_pb_pop_valid; // @[Scheduler.scala 53:21]
  wire [1:0] sinkA_io_pb_pop_bits_index; // @[Scheduler.scala 53:21]
  wire [255:0] sinkA_io_pb_beat_data; // @[Scheduler.scala 53:21]
  wire [7:0] sinkA_io_pb_beat_mask; // @[Scheduler.scala 53:21]
  wire  sinkA_io_pb_pop2_ready; // @[Scheduler.scala 53:21]
  wire  sinkA_io_pb_pop2_valid; // @[Scheduler.scala 53:21]
  wire [1:0] sinkA_io_pb_pop2_bits_index; // @[Scheduler.scala 53:21]
  wire [255:0] sinkA_io_pb_beat2_data; // @[Scheduler.scala 53:21]
  wire [7:0] sinkA_io_pb_beat2_mask; // @[Scheduler.scala 53:21]
  wire  sinkD_clock; // @[Scheduler.scala 54:21]
  wire  sinkD_reset; // @[Scheduler.scala 54:21]
  wire  sinkD_io_resp_valid; // @[Scheduler.scala 54:21]
  wire [2:0] sinkD_io_resp_bits_opcode; // @[Scheduler.scala 54:21]
  wire [3:0] sinkD_io_resp_bits_source; // @[Scheduler.scala 54:21]
  wire [255:0] sinkD_io_resp_bits_data; // @[Scheduler.scala 54:21]
  wire  sinkD_io_d_ready; // @[Scheduler.scala 54:21]
  wire  sinkD_io_d_valid; // @[Scheduler.scala 54:21]
  wire [2:0] sinkD_io_d_bits_opcode; // @[Scheduler.scala 54:21]
  wire [3:0] sinkD_io_d_bits_source; // @[Scheduler.scala 54:21]
  wire [255:0] sinkD_io_d_bits_data; // @[Scheduler.scala 54:21]
  wire [3:0] sinkD_io_source; // @[Scheduler.scala 54:21]
  wire [1:0] sinkD_io_way; // @[Scheduler.scala 54:21]
  wire  sinkD_io_set; // @[Scheduler.scala 54:21]
  wire [2:0] sinkD_io_opcode; // @[Scheduler.scala 54:21]
  wire [1:0] sinkD_io_put; // @[Scheduler.scala 54:21]
  wire  sinkD_io_bs_adr_valid; // @[Scheduler.scala 54:21]
  wire [1:0] sinkD_io_bs_adr_bits_way; // @[Scheduler.scala 54:21]
  wire  sinkD_io_bs_adr_bits_set; // @[Scheduler.scala 54:21]
  wire [255:0] sinkD_io_bs_dat_data; // @[Scheduler.scala 54:21]
  wire  sinkD_io_pb_pop_valid; // @[Scheduler.scala 54:21]
  wire [1:0] sinkD_io_pb_pop_bits_index; // @[Scheduler.scala 54:21]
  wire [255:0] sinkD_io_pb_beat_data; // @[Scheduler.scala 54:21]
  wire [7:0] sinkD_io_pb_beat_mask; // @[Scheduler.scala 54:21]
  wire  directory_clock; // @[Scheduler.scala 89:25]
  wire  directory_reset; // @[Scheduler.scala 89:25]
  wire  directory_io_write_ready; // @[Scheduler.scala 89:25]
  wire  directory_io_write_valid; // @[Scheduler.scala 89:25]
  wire [1:0] directory_io_write_bits_way; // @[Scheduler.scala 89:25]
  wire [25:0] directory_io_write_bits_data_tag; // @[Scheduler.scala 89:25]
  wire  directory_io_write_bits_data_valid; // @[Scheduler.scala 89:25]
  wire  directory_io_write_bits_set; // @[Scheduler.scala 89:25]
  wire  directory_io_read_ready; // @[Scheduler.scala 89:25]
  wire  directory_io_read_valid; // @[Scheduler.scala 89:25]
  wire [2:0] directory_io_read_bits_opcode; // @[Scheduler.scala 89:25]
  wire [3:0] directory_io_read_bits_source; // @[Scheduler.scala 89:25]
  wire [25:0] directory_io_read_bits_tag; // @[Scheduler.scala 89:25]
  wire [4:0] directory_io_read_bits_offset; // @[Scheduler.scala 89:25]
  wire [1:0] directory_io_read_bits_put; // @[Scheduler.scala 89:25]
  wire [255:0] directory_io_read_bits_data; // @[Scheduler.scala 89:25]
  wire [7:0] directory_io_read_bits_mask; // @[Scheduler.scala 89:25]
  wire  directory_io_read_bits_set; // @[Scheduler.scala 89:25]
  wire  directory_io_result_valid; // @[Scheduler.scala 89:25]
  wire [2:0] directory_io_result_bits_opcode; // @[Scheduler.scala 89:25]
  wire [3:0] directory_io_result_bits_source; // @[Scheduler.scala 89:25]
  wire [25:0] directory_io_result_bits_tag; // @[Scheduler.scala 89:25]
  wire [4:0] directory_io_result_bits_offset; // @[Scheduler.scala 89:25]
  wire [1:0] directory_io_result_bits_put; // @[Scheduler.scala 89:25]
  wire [255:0] directory_io_result_bits_data; // @[Scheduler.scala 89:25]
  wire [7:0] directory_io_result_bits_mask; // @[Scheduler.scala 89:25]
  wire  directory_io_result_bits_set; // @[Scheduler.scala 89:25]
  wire  directory_io_result_bits_hit; // @[Scheduler.scala 89:25]
  wire [1:0] directory_io_result_bits_way; // @[Scheduler.scala 89:25]
  wire  bankedStore_clock; // @[Scheduler.scala 91:27]
  wire  bankedStore_reset; // @[Scheduler.scala 91:27]
  wire  bankedStore_io_sinkD_adr_valid; // @[Scheduler.scala 91:27]
  wire [1:0] bankedStore_io_sinkD_adr_bits_way; // @[Scheduler.scala 91:27]
  wire  bankedStore_io_sinkD_adr_bits_set; // @[Scheduler.scala 91:27]
  wire [255:0] bankedStore_io_sinkD_dat_data; // @[Scheduler.scala 91:27]
  wire  bankedStore_io_sourceD_radr_valid; // @[Scheduler.scala 91:27]
  wire [1:0] bankedStore_io_sourceD_radr_bits_way; // @[Scheduler.scala 91:27]
  wire  bankedStore_io_sourceD_radr_bits_set; // @[Scheduler.scala 91:27]
  wire [7:0] bankedStore_io_sourceD_radr_bits_mask; // @[Scheduler.scala 91:27]
  wire [255:0] bankedStore_io_sourceD_rdat_data; // @[Scheduler.scala 91:27]
  wire  bankedStore_io_sourceD_wadr_valid; // @[Scheduler.scala 91:27]
  wire [1:0] bankedStore_io_sourceD_wadr_bits_way; // @[Scheduler.scala 91:27]
  wire  bankedStore_io_sourceD_wadr_bits_set; // @[Scheduler.scala 91:27]
  wire [7:0] bankedStore_io_sourceD_wadr_bits_mask; // @[Scheduler.scala 91:27]
  wire [255:0] bankedStore_io_sourceD_wdat_data; // @[Scheduler.scala 91:27]
  wire  requests_clock; // @[Scheduler.scala 94:24]
  wire  requests_reset; // @[Scheduler.scala 94:24]
  wire  requests_io_push_ready; // @[Scheduler.scala 94:24]
  wire  requests_io_push_valid; // @[Scheduler.scala 94:24]
  wire [1:0] requests_io_push_bits_index; // @[Scheduler.scala 94:24]
  wire [3:0] requests_io_push_bits_data; // @[Scheduler.scala 94:24]
  wire [3:0] requests_io_valid; // @[Scheduler.scala 94:24]
  wire  requests_io_pop_valid; // @[Scheduler.scala 94:24]
  wire [1:0] requests_io_pop_bits; // @[Scheduler.scala 94:24]
  wire [3:0] requests_io_data; // @[Scheduler.scala 94:24]
  wire  mshrs_0_clock; // @[Scheduler.scala 96:46]
  wire  mshrs_0_reset; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_allocate_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_0_io_allocate_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_0_io_allocate_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_0_io_allocate_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_allocate_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_0_io_allocate_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_0_io_allocate_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_allocate_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_allocate_bits_way; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_0_io_status_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_0_io_status_tag; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_status_put; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_status_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_status_way; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_valid; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_a_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_a_valid; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_0_io_schedule_a_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_0_io_schedule_a_bits_offset; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_0_io_schedule_a_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_a_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_d_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_0_io_schedule_d_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_0_io_schedule_d_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_0_io_schedule_d_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_schedule_d_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_0_io_schedule_d_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_0_io_schedule_d_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_d_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_schedule_d_bits_way; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_dir_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_dir_valid; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_0_io_schedule_dir_bits_way; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_0_io_schedule_dir_bits_data_tag; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_schedule_dir_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_0_io_sinkd_valid; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_0_io_sinkd_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_1_clock; // @[Scheduler.scala 96:46]
  wire  mshrs_1_reset; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_allocate_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_1_io_allocate_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_1_io_allocate_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_1_io_allocate_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_allocate_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_1_io_allocate_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_1_io_allocate_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_allocate_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_allocate_bits_way; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_1_io_status_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_1_io_status_tag; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_status_put; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_status_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_status_way; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_valid; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_a_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_a_valid; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_1_io_schedule_a_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_1_io_schedule_a_bits_offset; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_1_io_schedule_a_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_a_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_d_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_1_io_schedule_d_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_1_io_schedule_d_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_1_io_schedule_d_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_schedule_d_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_1_io_schedule_d_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_1_io_schedule_d_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_d_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_schedule_d_bits_way; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_dir_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_dir_valid; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_1_io_schedule_dir_bits_way; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_1_io_schedule_dir_bits_data_tag; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_schedule_dir_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_1_io_sinkd_valid; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_1_io_sinkd_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_2_clock; // @[Scheduler.scala 96:46]
  wire  mshrs_2_reset; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_allocate_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_2_io_allocate_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_2_io_allocate_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_2_io_allocate_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_allocate_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_2_io_allocate_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_2_io_allocate_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_allocate_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_allocate_bits_way; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_2_io_status_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_2_io_status_tag; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_status_put; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_status_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_status_way; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_valid; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_a_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_a_valid; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_2_io_schedule_a_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_2_io_schedule_a_bits_offset; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_2_io_schedule_a_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_a_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_d_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_2_io_schedule_d_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_2_io_schedule_d_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_2_io_schedule_d_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_schedule_d_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_2_io_schedule_d_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_2_io_schedule_d_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_d_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_schedule_d_bits_way; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_dir_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_dir_valid; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_2_io_schedule_dir_bits_way; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_2_io_schedule_dir_bits_data_tag; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_schedule_dir_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_2_io_sinkd_valid; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_2_io_sinkd_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_3_clock; // @[Scheduler.scala 96:46]
  wire  mshrs_3_reset; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_allocate_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_3_io_allocate_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_3_io_allocate_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_3_io_allocate_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_allocate_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_3_io_allocate_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_3_io_allocate_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_allocate_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_allocate_bits_way; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_3_io_status_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_3_io_status_tag; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_status_put; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_status_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_status_way; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_valid; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_a_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_a_valid; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_3_io_schedule_a_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_3_io_schedule_a_bits_offset; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_3_io_schedule_a_bits_data; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_a_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_d_valid; // @[Scheduler.scala 96:46]
  wire [2:0] mshrs_3_io_schedule_d_bits_opcode; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_3_io_schedule_d_bits_tag; // @[Scheduler.scala 96:46]
  wire [4:0] mshrs_3_io_schedule_d_bits_offset; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_schedule_d_bits_put; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_3_io_schedule_d_bits_data; // @[Scheduler.scala 96:46]
  wire [7:0] mshrs_3_io_schedule_d_bits_mask; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_d_bits_set; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_schedule_d_bits_way; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_dir_ready; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_dir_valid; // @[Scheduler.scala 96:46]
  wire [1:0] mshrs_3_io_schedule_dir_bits_way; // @[Scheduler.scala 96:46]
  wire [25:0] mshrs_3_io_schedule_dir_bits_data_tag; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_schedule_dir_bits_set; // @[Scheduler.scala 96:46]
  wire  mshrs_3_io_sinkd_valid; // @[Scheduler.scala 96:46]
  wire [255:0] mshrs_3_io_sinkd_bits_data; // @[Scheduler.scala 96:46]
  wire  write_buffer_clock; // @[Scheduler.scala 140:27]
  wire  write_buffer_reset; // @[Scheduler.scala 140:27]
  wire  write_buffer_io_enq_ready; // @[Scheduler.scala 140:27]
  wire  write_buffer_io_enq_valid; // @[Scheduler.scala 140:27]
  wire [3:0] write_buffer_io_enq_bits_source; // @[Scheduler.scala 140:27]
  wire [25:0] write_buffer_io_enq_bits_tag; // @[Scheduler.scala 140:27]
  wire [4:0] write_buffer_io_enq_bits_offset; // @[Scheduler.scala 140:27]
  wire [255:0] write_buffer_io_enq_bits_data; // @[Scheduler.scala 140:27]
  wire [7:0] write_buffer_io_enq_bits_mask; // @[Scheduler.scala 140:27]
  wire  write_buffer_io_enq_bits_set; // @[Scheduler.scala 140:27]
  wire  write_buffer_io_deq_ready; // @[Scheduler.scala 140:27]
  wire  write_buffer_io_deq_valid; // @[Scheduler.scala 140:27]
  wire [2:0] write_buffer_io_deq_bits_opcode; // @[Scheduler.scala 140:27]
  wire [3:0] write_buffer_io_deq_bits_source; // @[Scheduler.scala 140:27]
  wire [25:0] write_buffer_io_deq_bits_tag; // @[Scheduler.scala 140:27]
  wire [4:0] write_buffer_io_deq_bits_offset; // @[Scheduler.scala 140:27]
  wire [255:0] write_buffer_io_deq_bits_data; // @[Scheduler.scala 140:27]
  wire [7:0] write_buffer_io_deq_bits_mask; // @[Scheduler.scala 140:27]
  wire  write_buffer_io_deq_bits_set; // @[Scheduler.scala 140:27]
  wire  dir_result_buffer_clock; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_reset; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_enq_ready; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_enq_valid; // @[Scheduler.scala 211:31]
  wire [2:0] dir_result_buffer_io_enq_bits_opcode; // @[Scheduler.scala 211:31]
  wire [3:0] dir_result_buffer_io_enq_bits_source; // @[Scheduler.scala 211:31]
  wire [25:0] dir_result_buffer_io_enq_bits_tag; // @[Scheduler.scala 211:31]
  wire [4:0] dir_result_buffer_io_enq_bits_offset; // @[Scheduler.scala 211:31]
  wire [1:0] dir_result_buffer_io_enq_bits_put; // @[Scheduler.scala 211:31]
  wire [255:0] dir_result_buffer_io_enq_bits_data; // @[Scheduler.scala 211:31]
  wire [7:0] dir_result_buffer_io_enq_bits_mask; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_enq_bits_set; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_enq_bits_hit; // @[Scheduler.scala 211:31]
  wire [1:0] dir_result_buffer_io_enq_bits_way; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_deq_ready; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_deq_valid; // @[Scheduler.scala 211:31]
  wire [2:0] dir_result_buffer_io_deq_bits_opcode; // @[Scheduler.scala 211:31]
  wire [3:0] dir_result_buffer_io_deq_bits_source; // @[Scheduler.scala 211:31]
  wire [25:0] dir_result_buffer_io_deq_bits_tag; // @[Scheduler.scala 211:31]
  wire [4:0] dir_result_buffer_io_deq_bits_offset; // @[Scheduler.scala 211:31]
  wire [1:0] dir_result_buffer_io_deq_bits_put; // @[Scheduler.scala 211:31]
  wire [255:0] dir_result_buffer_io_deq_bits_data; // @[Scheduler.scala 211:31]
  wire [7:0] dir_result_buffer_io_deq_bits_mask; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_deq_bits_set; // @[Scheduler.scala 211:31]
  wire  dir_result_buffer_io_deq_bits_hit; // @[Scheduler.scala 211:31]
  wire [1:0] dir_result_buffer_io_deq_bits_way; // @[Scheduler.scala 211:31]
  wire [1:0] _sinkD_io_way_WIRE_0 = mshrs_0_io_status_way; // @[Scheduler.scala 100:{28,28}]
  wire [1:0] _sinkD_io_way_WIRE_1 = mshrs_1_io_status_way; // @[Scheduler.scala 100:{28,28}]
  wire [1:0] _GEN_1 = 2'h1 == sinkD_io_source[1:0] ? _sinkD_io_way_WIRE_1 : _sinkD_io_way_WIRE_0; // @[Scheduler.scala 100:{18,18}]
  wire [1:0] _sinkD_io_way_WIRE_2 = mshrs_2_io_status_way; // @[Scheduler.scala 100:{28,28}]
  wire [1:0] _GEN_2 = 2'h2 == sinkD_io_source[1:0] ? _sinkD_io_way_WIRE_2 : _GEN_1; // @[Scheduler.scala 100:{18,18}]
  wire [1:0] _sinkD_io_way_WIRE_3 = mshrs_3_io_status_way; // @[Scheduler.scala 100:{28,28}]
  wire  _GEN_5 = 2'h1 == sinkD_io_source[1:0] ? mshrs_1_io_status_set : mshrs_0_io_status_set; // @[Scheduler.scala 101:{18,18}]
  wire  _GEN_6 = 2'h2 == sinkD_io_source[1:0] ? mshrs_2_io_status_set : _GEN_5; // @[Scheduler.scala 101:{18,18}]
  wire [2:0] _sinkD_io_opcode_WIRE_0 = mshrs_0_io_status_opcode; // @[Scheduler.scala 102:{28,28}]
  wire [2:0] _sinkD_io_opcode_WIRE_1 = mshrs_1_io_status_opcode; // @[Scheduler.scala 102:{28,28}]
  wire [2:0] _GEN_9 = 2'h1 == sinkD_io_source[1:0] ? _sinkD_io_opcode_WIRE_1 : _sinkD_io_opcode_WIRE_0; // @[Scheduler.scala 102:{18,18}]
  wire [2:0] _sinkD_io_opcode_WIRE_2 = mshrs_2_io_status_opcode; // @[Scheduler.scala 102:{28,28}]
  wire [2:0] _GEN_10 = 2'h2 == sinkD_io_source[1:0] ? _sinkD_io_opcode_WIRE_2 : _GEN_9; // @[Scheduler.scala 102:{18,18}]
  wire [2:0] _sinkD_io_opcode_WIRE_3 = mshrs_3_io_status_opcode; // @[Scheduler.scala 102:{28,28}]
  wire [1:0] _sinkD_io_put_WIRE_0 = mshrs_0_io_status_put; // @[Scheduler.scala 103:{28,28}]
  wire [1:0] _sinkD_io_put_WIRE_1 = mshrs_1_io_status_put; // @[Scheduler.scala 103:{28,28}]
  wire [1:0] _GEN_13 = 2'h1 == sinkD_io_source[1:0] ? _sinkD_io_put_WIRE_1 : _sinkD_io_put_WIRE_0; // @[Scheduler.scala 103:{18,18}]
  wire [1:0] _sinkD_io_put_WIRE_2 = mshrs_2_io_status_put; // @[Scheduler.scala 103:{28,28}]
  wire [1:0] _GEN_14 = 2'h2 == sinkD_io_source[1:0] ? _sinkD_io_put_WIRE_2 : _GEN_13; // @[Scheduler.scala 103:{18,18}]
  wire [1:0] _sinkD_io_put_WIRE_3 = mshrs_3_io_status_put; // @[Scheduler.scala 103:{28,28}]
  wire  _mshr_request_T_1 = sourceD_io_req_ready & mshrs_0_io_schedule_d_valid; // @[Scheduler.scala 107:29]
  wire  _mshr_request_T_2 = sourceA_io_req_ready & mshrs_0_io_schedule_a_valid | _mshr_request_T_1; // @[Scheduler.scala 106:54]
  wire  _mshr_request_T_3 = mshrs_0_io_schedule_dir_valid & directory_io_write_ready; // @[Scheduler.scala 109:31]
  wire  _mshr_request_T_4 = _mshr_request_T_2 | _mshr_request_T_3; // @[Scheduler.scala 107:54]
  wire  _mshr_request_T_6 = sourceD_io_req_ready & mshrs_1_io_schedule_d_valid; // @[Scheduler.scala 107:29]
  wire  _mshr_request_T_7 = sourceA_io_req_ready & mshrs_1_io_schedule_a_valid | _mshr_request_T_6; // @[Scheduler.scala 106:54]
  wire  _mshr_request_T_8 = mshrs_1_io_schedule_dir_valid & directory_io_write_ready; // @[Scheduler.scala 109:31]
  wire  _mshr_request_T_9 = _mshr_request_T_7 | _mshr_request_T_8; // @[Scheduler.scala 107:54]
  wire  _mshr_request_T_11 = sourceD_io_req_ready & mshrs_2_io_schedule_d_valid; // @[Scheduler.scala 107:29]
  wire  _mshr_request_T_12 = sourceA_io_req_ready & mshrs_2_io_schedule_a_valid | _mshr_request_T_11; // @[Scheduler.scala 106:54]
  wire  _mshr_request_T_13 = mshrs_2_io_schedule_dir_valid & directory_io_write_ready; // @[Scheduler.scala 109:31]
  wire  _mshr_request_T_14 = _mshr_request_T_12 | _mshr_request_T_13; // @[Scheduler.scala 107:54]
  wire  _mshr_request_T_16 = sourceD_io_req_ready & mshrs_3_io_schedule_d_valid; // @[Scheduler.scala 107:29]
  wire  _mshr_request_T_17 = sourceA_io_req_ready & mshrs_3_io_schedule_a_valid | _mshr_request_T_16; // @[Scheduler.scala 106:54]
  wire  _mshr_request_T_18 = mshrs_3_io_schedule_dir_valid & directory_io_write_ready; // @[Scheduler.scala 109:31]
  wire  _mshr_request_T_19 = _mshr_request_T_17 | _mshr_request_T_18; // @[Scheduler.scala 107:54]
  wire [3:0] mshr_request = {_mshr_request_T_19,_mshr_request_T_14,_mshr_request_T_9,_mshr_request_T_4}; // @[Cat.scala 31:58]
  reg [3:0] robin_filter; // @[Scheduler.scala 113:29]
  wire [3:0] _robin_request_T = mshr_request & robin_filter; // @[Scheduler.scala 114:54]
  wire [7:0] robin_request = {_mshr_request_T_19,_mshr_request_T_14,_mshr_request_T_9,_mshr_request_T_4,_robin_request_T
    }; // @[Cat.scala 31:58]
  wire [8:0] _mshr_selectOH2_T = {robin_request, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _mshr_selectOH2_T_2 = robin_request | _mshr_selectOH2_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _mshr_selectOH2_T_3 = {_mshr_selectOH2_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _mshr_selectOH2_T_5 = _mshr_selectOH2_T_2 | _mshr_selectOH2_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _mshr_selectOH2_T_6 = {_mshr_selectOH2_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _mshr_selectOH2_T_8 = _mshr_selectOH2_T_5 | _mshr_selectOH2_T_6[7:0]; // @[package.scala 244:43]
  wire [8:0] _mshr_selectOH2_T_10 = {_mshr_selectOH2_T_8, 1'h0}; // @[Scheduler.scala 115:49]
  wire [8:0] _mshr_selectOH2_T_11 = ~_mshr_selectOH2_T_10; // @[Scheduler.scala 115:25]
  wire [8:0] _GEN_65 = {{1'd0}, robin_request}; // @[Scheduler.scala 115:65]
  wire [8:0] mshr_selectOH2 = _mshr_selectOH2_T_11 & _GEN_65; // @[Scheduler.scala 115:65]
  wire [3:0] mshr_selectOH = mshr_selectOH2[7:4] | mshr_selectOH2[3:0]; // @[Scheduler.scala 116:70]
  wire [1:0] mshr_select_hi = mshr_selectOH[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] mshr_select_lo = mshr_selectOH[1:0]; // @[OneHot.scala 31:18]
  wire  _mshr_select_T = |mshr_select_hi; // @[OneHot.scala 32:14]
  wire [1:0] _mshr_select_T_1 = mshr_select_hi | mshr_select_lo; // @[OneHot.scala 32:28]
  wire [1:0] mshr_select = {_mshr_select_T,_mshr_select_T_1[1]}; // @[Cat.scala 31:58]
  wire [25:0] _schedule_T_18 = mshr_selectOH[0] ? mshrs_0_io_schedule_dir_bits_data_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_19 = mshr_selectOH[1] ? mshrs_1_io_schedule_dir_bits_data_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_20 = mshr_selectOH[2] ? mshrs_2_io_schedule_dir_bits_data_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_21 = mshr_selectOH[3] ? mshrs_3_io_schedule_dir_bits_data_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_22 = _schedule_T_18 | _schedule_T_19; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_23 = _schedule_T_22 | _schedule_T_20; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_25 = mshr_selectOH[0] ? mshrs_0_io_schedule_dir_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_26 = mshr_selectOH[1] ? mshrs_1_io_schedule_dir_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_27 = mshr_selectOH[2] ? mshrs_2_io_schedule_dir_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_28 = mshr_selectOH[3] ? mshrs_3_io_schedule_dir_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_29 = _schedule_T_25 | _schedule_T_26; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_30 = _schedule_T_29 | _schedule_T_27; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_46 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_47 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_48 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_49 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_way : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_50 = _schedule_T_46 | _schedule_T_47; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_51 = _schedule_T_50 | _schedule_T_48; // @[Mux.scala 27:73]
  wire [1:0] schedule_d_bits_way = _schedule_T_51 | _schedule_T_49; // @[Mux.scala 27:73]
  wire  schedule_d_bits_set = mshr_selectOH[0] & mshrs_0_io_schedule_d_bits_set | mshr_selectOH[1] &
    mshrs_1_io_schedule_d_bits_set | mshr_selectOH[2] & mshrs_2_io_schedule_d_bits_set | mshr_selectOH[3] &
    mshrs_3_io_schedule_d_bits_set; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_67 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_68 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_69 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_70 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_71 = _schedule_T_67 | _schedule_T_68; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_72 = _schedule_T_71 | _schedule_T_69; // @[Mux.scala 27:73]
  wire [7:0] schedule_d_bits_mask = _schedule_T_72 | _schedule_T_70; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_74 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_75 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_76 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_77 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_78 = _schedule_T_74 | _schedule_T_75; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_79 = _schedule_T_78 | _schedule_T_76; // @[Mux.scala 27:73]
  wire [255:0] schedule_d_bits_data = _schedule_T_79 | _schedule_T_77; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_81 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_put : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_82 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_put : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_83 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_put : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_84 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_put : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_85 = _schedule_T_81 | _schedule_T_82; // @[Mux.scala 27:73]
  wire [1:0] _schedule_T_86 = _schedule_T_85 | _schedule_T_83; // @[Mux.scala 27:73]
  wire [1:0] schedule_d_bits_put = _schedule_T_86 | _schedule_T_84; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_88 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_89 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_90 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_91 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_92 = _schedule_T_88 | _schedule_T_89; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_93 = _schedule_T_92 | _schedule_T_90; // @[Mux.scala 27:73]
  wire [4:0] schedule_d_bits_offset = _schedule_T_93 | _schedule_T_91; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_95 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_96 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_97 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_98 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_99 = _schedule_T_95 | _schedule_T_96; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_100 = _schedule_T_99 | _schedule_T_97; // @[Mux.scala 27:73]
  wire [25:0] schedule_d_bits_tag = _schedule_T_100 | _schedule_T_98; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_116 = mshr_selectOH[0] ? mshrs_0_io_schedule_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_117 = mshr_selectOH[1] ? mshrs_1_io_schedule_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_118 = mshr_selectOH[2] ? mshrs_2_io_schedule_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_119 = mshr_selectOH[3] ? mshrs_3_io_schedule_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_120 = _schedule_T_116 | _schedule_T_117; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_121 = _schedule_T_120 | _schedule_T_118; // @[Mux.scala 27:73]
  wire [2:0] schedule_d_bits_opcode = _schedule_T_121 | _schedule_T_119; // @[Mux.scala 27:73]
  wire  schedule_d_valid = mshr_selectOH[0] & mshrs_0_io_schedule_d_valid | mshr_selectOH[1] &
    mshrs_1_io_schedule_d_valid | mshr_selectOH[2] & mshrs_2_io_schedule_d_valid | mshr_selectOH[3] &
    mshrs_3_io_schedule_d_valid; // @[Mux.scala 27:73]
  wire  schedule_a_bits_set = mshr_selectOH[0] & mshrs_0_io_schedule_a_bits_set | mshr_selectOH[1] &
    mshrs_1_io_schedule_a_bits_set | mshr_selectOH[2] & mshrs_2_io_schedule_a_bits_set | mshr_selectOH[3] &
    mshrs_3_io_schedule_a_bits_set; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_144 = mshr_selectOH[0] ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_145 = mshr_selectOH[1] ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_146 = mshr_selectOH[2] ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_147 = mshr_selectOH[3] ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_148 = _schedule_T_144 | _schedule_T_145; // @[Mux.scala 27:73]
  wire [7:0] _schedule_T_149 = _schedule_T_148 | _schedule_T_146; // @[Mux.scala 27:73]
  wire [7:0] schedule_a_bits_mask = _schedule_T_149 | _schedule_T_147; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_151 = mshr_selectOH[0] ? mshrs_0_io_schedule_a_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_152 = mshr_selectOH[1] ? mshrs_1_io_schedule_a_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_153 = mshr_selectOH[2] ? mshrs_2_io_schedule_a_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_154 = mshr_selectOH[3] ? mshrs_3_io_schedule_a_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_155 = _schedule_T_151 | _schedule_T_152; // @[Mux.scala 27:73]
  wire [255:0] _schedule_T_156 = _schedule_T_155 | _schedule_T_153; // @[Mux.scala 27:73]
  wire [255:0] schedule_a_bits_data = _schedule_T_156 | _schedule_T_154; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_165 = mshr_selectOH[0] ? mshrs_0_io_schedule_a_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_166 = mshr_selectOH[1] ? mshrs_1_io_schedule_a_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_167 = mshr_selectOH[2] ? mshrs_2_io_schedule_a_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_168 = mshr_selectOH[3] ? mshrs_3_io_schedule_a_bits_offset : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_169 = _schedule_T_165 | _schedule_T_166; // @[Mux.scala 27:73]
  wire [4:0] _schedule_T_170 = _schedule_T_169 | _schedule_T_167; // @[Mux.scala 27:73]
  wire [4:0] schedule_a_bits_offset = _schedule_T_170 | _schedule_T_168; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_172 = mshr_selectOH[0] ? mshrs_0_io_schedule_a_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_173 = mshr_selectOH[1] ? mshrs_1_io_schedule_a_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_174 = mshr_selectOH[2] ? mshrs_2_io_schedule_a_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_175 = mshr_selectOH[3] ? mshrs_3_io_schedule_a_bits_tag : 26'h0; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_176 = _schedule_T_172 | _schedule_T_173; // @[Mux.scala 27:73]
  wire [25:0] _schedule_T_177 = _schedule_T_176 | _schedule_T_174; // @[Mux.scala 27:73]
  wire [25:0] schedule_a_bits_tag = _schedule_T_177 | _schedule_T_175; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_193 = mshr_selectOH[0] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_194 = mshr_selectOH[1] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_195 = mshr_selectOH[2] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_196 = mshr_selectOH[3] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_197 = _schedule_T_193 | _schedule_T_194; // @[Mux.scala 27:73]
  wire [2:0] _schedule_T_198 = _schedule_T_197 | _schedule_T_195; // @[Mux.scala 27:73]
  wire [2:0] schedule_a_bits_opcode = _schedule_T_198 | _schedule_T_196; // @[Mux.scala 27:73]
  wire  schedule_a_valid = mshr_selectOH[0] & mshrs_0_io_schedule_a_valid | mshr_selectOH[1] &
    mshrs_1_io_schedule_a_valid | mshr_selectOH[2] & mshrs_2_io_schedule_a_valid | mshr_selectOH[3] &
    mshrs_3_io_schedule_a_valid; // @[Mux.scala 27:73]
  wire [3:0] _GEN_66 = {{1'd0}, mshr_selectOH[3:1]}; // @[package.scala 253:43]
  wire [3:0] _robin_filter_T_1 = mshr_selectOH | _GEN_66; // @[package.scala 253:43]
  wire [3:0] _GEN_67 = {{2'd0}, _robin_filter_T_1[3:2]}; // @[package.scala 253:43]
  wire [3:0] _robin_filter_T_3 = _robin_filter_T_1 | _GEN_67; // @[package.scala 253:43]
  wire [3:0] _robin_filter_T_5 = ~_robin_filter_T_3; // @[Scheduler.scala 124:47]
  wire  _mshrs_0_io_schedule_a_ready_T = mshr_select == 2'h0; // @[Scheduler.scala 132:65]
  wire  _mshrs_1_io_schedule_a_ready_T = mshr_select == 2'h1; // @[Scheduler.scala 132:65]
  wire  _mshrs_2_io_schedule_a_ready_T = mshr_select == 2'h2; // @[Scheduler.scala 132:65]
  wire  _mshrs_3_io_schedule_a_ready_T = mshr_select == 2'h3; // @[Scheduler.scala 132:65]
  wire [3:0] schedule_a_bits_source = {{2'd0}, mshr_select}; // @[Mux.scala 27:73 Scheduler.scala 127:26]
  wire  _tagMatches_T_3 = ~directory_io_result_bits_hit; // @[Scheduler.scala 176:140]
  wire  _tagMatches_T_4 = requests_io_valid[0] & mshrs_0_io_status_tag == directory_io_result_bits_tag & ~
    directory_io_result_bits_hit; // @[Scheduler.scala 176:136]
  wire  _tagMatches_T_9 = requests_io_valid[1] & mshrs_1_io_status_tag == directory_io_result_bits_tag & ~
    directory_io_result_bits_hit; // @[Scheduler.scala 176:136]
  wire  _tagMatches_T_14 = requests_io_valid[2] & mshrs_2_io_status_tag == directory_io_result_bits_tag & ~
    directory_io_result_bits_hit; // @[Scheduler.scala 176:136]
  wire  _tagMatches_T_19 = requests_io_valid[3] & mshrs_3_io_status_tag == directory_io_result_bits_tag & ~
    directory_io_result_bits_hit; // @[Scheduler.scala 176:136]
  wire [3:0] tagMatches = {_tagMatches_T_19,_tagMatches_T_14,_tagMatches_T_9,_tagMatches_T_4}; // @[Cat.scala 31:58]
  wire  alloc = ~(|tagMatches); // @[Scheduler.scala 177:15]
  wire [3:0] _mshr_free_T = ~requests_io_valid; // @[Scheduler.scala 180:20]
  wire  mshr_free = |_mshr_free_T; // @[Scheduler.scala 180:45]
  wire [4:0] _mshr_insertOH_init_T_1 = {_mshr_free_T, 1'h0}; // @[package.scala 244:48]
  wire [3:0] _mshr_insertOH_init_T_3 = _mshr_free_T | _mshr_insertOH_init_T_1[3:0]; // @[package.scala 244:43]
  wire [5:0] _mshr_insertOH_init_T_4 = {_mshr_insertOH_init_T_3, 2'h0}; // @[package.scala 244:48]
  wire [3:0] _mshr_insertOH_init_T_6 = _mshr_insertOH_init_T_3 | _mshr_insertOH_init_T_4[3:0]; // @[package.scala 244:43]
  wire [4:0] _mshr_insertOH_init_T_8 = {_mshr_insertOH_init_T_6, 1'h0}; // @[Scheduler.scala 184:63]
  wire [4:0] _mshr_insertOH_init_T_9 = ~_mshr_insertOH_init_T_8; // @[Scheduler.scala 184:29]
  wire [4:0] _GEN_68 = {{1'd0}, _mshr_free_T}; // @[Scheduler.scala 184:79]
  wire [4:0] mshr_insertOH = _mshr_insertOH_init_T_9 & _GEN_68; // @[Scheduler.scala 184:79]
  wire [4:0] _requests_io_push_bits_index_T = alloc ? mshr_insertOH : {{1'd0}, tagMatches}; // @[Scheduler.scala 197:46]
  wire  requests_io_push_bits_index_hi = _requests_io_push_bits_index_T[4]; // @[OneHot.scala 30:18]
  wire [3:0] requests_io_push_bits_index_lo = _requests_io_push_bits_index_T[3:0]; // @[OneHot.scala 31:18]
  wire  _requests_io_push_bits_index_T_1 = |requests_io_push_bits_index_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_69 = {{3'd0}, requests_io_push_bits_index_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _requests_io_push_bits_index_T_2 = _GEN_69 | requests_io_push_bits_index_lo; // @[OneHot.scala 32:28]
  wire [1:0] requests_io_push_bits_index_hi_1 = _requests_io_push_bits_index_T_2[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] requests_io_push_bits_index_lo_1 = _requests_io_push_bits_index_T_2[1:0]; // @[OneHot.scala 31:18]
  wire  _requests_io_push_bits_index_T_3 = |requests_io_push_bits_index_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _requests_io_push_bits_index_T_4 = requests_io_push_bits_index_hi_1 | requests_io_push_bits_index_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] _requests_io_push_bits_index_T_7 = {_requests_io_push_bits_index_T_1,_requests_io_push_bits_index_T_3,
    _requests_io_push_bits_index_T_4[1]}; // @[Cat.scala 31:58]
  wire [3:0] _requests_io_pop_valid_T = requests_io_valid >> mshr_select; // @[Scheduler.scala 202:45]
  wire  _dir_result_buffer_io_deq_ready_T = ~schedule_d_valid; // @[Scheduler.scala 215:36]
  SourceA sourceA ( // @[Scheduler.scala 49:23]
    .io_req_ready(sourceA_io_req_ready),
    .io_req_valid(sourceA_io_req_valid),
    .io_req_bits_opcode(sourceA_io_req_bits_opcode),
    .io_req_bits_source(sourceA_io_req_bits_source),
    .io_req_bits_tag(sourceA_io_req_bits_tag),
    .io_req_bits_offset(sourceA_io_req_bits_offset),
    .io_req_bits_data(sourceA_io_req_bits_data),
    .io_req_bits_mask(sourceA_io_req_bits_mask),
    .io_req_bits_set(sourceA_io_req_bits_set),
    .io_a_ready(sourceA_io_a_ready),
    .io_a_valid(sourceA_io_a_valid),
    .io_a_bits_opcode(sourceA_io_a_bits_opcode),
    .io_a_bits_source(sourceA_io_a_bits_source),
    .io_a_bits_address(sourceA_io_a_bits_address),
    .io_a_bits_mask(sourceA_io_a_bits_mask),
    .io_a_bits_data(sourceA_io_a_bits_data)
  );
  SourceD sourceD ( // @[Scheduler.scala 51:23]
    .clock(sourceD_clock),
    .reset(sourceD_reset),
    .io_req_ready(sourceD_io_req_ready),
    .io_req_valid(sourceD_io_req_valid),
    .io_req_bits_opcode(sourceD_io_req_bits_opcode),
    .io_req_bits_source(sourceD_io_req_bits_source),
    .io_req_bits_tag(sourceD_io_req_bits_tag),
    .io_req_bits_offset(sourceD_io_req_bits_offset),
    .io_req_bits_put(sourceD_io_req_bits_put),
    .io_req_bits_data(sourceD_io_req_bits_data),
    .io_req_bits_mask(sourceD_io_req_bits_mask),
    .io_req_bits_set(sourceD_io_req_bits_set),
    .io_req_bits_hit(sourceD_io_req_bits_hit),
    .io_req_bits_way(sourceD_io_req_bits_way),
    .io_req_bits_from_mem(sourceD_io_req_bits_from_mem),
    .io_d_ready(sourceD_io_d_ready),
    .io_d_valid(sourceD_io_d_valid),
    .io_d_bits_source(sourceD_io_d_bits_source),
    .io_d_bits_data(sourceD_io_d_bits_data),
    .io_d_bits_address(sourceD_io_d_bits_address),
    .io_pb_pop_valid(sourceD_io_pb_pop_valid),
    .io_pb_pop_bits_index(sourceD_io_pb_pop_bits_index),
    .io_pb_beat_data(sourceD_io_pb_beat_data),
    .io_pb_beat_mask(sourceD_io_pb_beat_mask),
    .io_bs_radr_valid(sourceD_io_bs_radr_valid),
    .io_bs_radr_bits_way(sourceD_io_bs_radr_bits_way),
    .io_bs_radr_bits_set(sourceD_io_bs_radr_bits_set),
    .io_bs_radr_bits_mask(sourceD_io_bs_radr_bits_mask),
    .io_bs_rdat_data(sourceD_io_bs_rdat_data),
    .io_bs_wadr_valid(sourceD_io_bs_wadr_valid),
    .io_bs_wadr_bits_way(sourceD_io_bs_wadr_bits_way),
    .io_bs_wadr_bits_set(sourceD_io_bs_wadr_bits_set),
    .io_bs_wadr_bits_mask(sourceD_io_bs_wadr_bits_mask),
    .io_bs_wdat_data(sourceD_io_bs_wdat_data),
    .io_a_ready(sourceD_io_a_ready),
    .io_a_valid(sourceD_io_a_valid),
    .io_a_bits_source(sourceD_io_a_bits_source),
    .io_a_bits_tag(sourceD_io_a_bits_tag),
    .io_a_bits_offset(sourceD_io_a_bits_offset),
    .io_a_bits_data(sourceD_io_a_bits_data),
    .io_a_bits_mask(sourceD_io_a_bits_mask),
    .io_a_bits_set(sourceD_io_a_bits_set)
  );
  SinkA sinkA ( // @[Scheduler.scala 53:21]
    .clock(sinkA_clock),
    .reset(sinkA_reset),
    .io_req_ready(sinkA_io_req_ready),
    .io_req_valid(sinkA_io_req_valid),
    .io_req_bits_opcode(sinkA_io_req_bits_opcode),
    .io_req_bits_source(sinkA_io_req_bits_source),
    .io_req_bits_tag(sinkA_io_req_bits_tag),
    .io_req_bits_offset(sinkA_io_req_bits_offset),
    .io_req_bits_put(sinkA_io_req_bits_put),
    .io_req_bits_data(sinkA_io_req_bits_data),
    .io_req_bits_mask(sinkA_io_req_bits_mask),
    .io_req_bits_set(sinkA_io_req_bits_set),
    .io_a_ready(sinkA_io_a_ready),
    .io_a_valid(sinkA_io_a_valid),
    .io_a_bits_opcode(sinkA_io_a_bits_opcode),
    .io_a_bits_source(sinkA_io_a_bits_source),
    .io_a_bits_address(sinkA_io_a_bits_address),
    .io_a_bits_mask(sinkA_io_a_bits_mask),
    .io_a_bits_data(sinkA_io_a_bits_data),
    .io_pb_pop_ready(sinkA_io_pb_pop_ready),
    .io_pb_pop_valid(sinkA_io_pb_pop_valid),
    .io_pb_pop_bits_index(sinkA_io_pb_pop_bits_index),
    .io_pb_beat_data(sinkA_io_pb_beat_data),
    .io_pb_beat_mask(sinkA_io_pb_beat_mask),
    .io_pb_pop2_ready(sinkA_io_pb_pop2_ready),
    .io_pb_pop2_valid(sinkA_io_pb_pop2_valid),
    .io_pb_pop2_bits_index(sinkA_io_pb_pop2_bits_index),
    .io_pb_beat2_data(sinkA_io_pb_beat2_data),
    .io_pb_beat2_mask(sinkA_io_pb_beat2_mask)
  );
  SinkD sinkD ( // @[Scheduler.scala 54:21]
    .clock(sinkD_clock),
    .reset(sinkD_reset),
    .io_resp_valid(sinkD_io_resp_valid),
    .io_resp_bits_opcode(sinkD_io_resp_bits_opcode),
    .io_resp_bits_source(sinkD_io_resp_bits_source),
    .io_resp_bits_data(sinkD_io_resp_bits_data),
    .io_d_ready(sinkD_io_d_ready),
    .io_d_valid(sinkD_io_d_valid),
    .io_d_bits_opcode(sinkD_io_d_bits_opcode),
    .io_d_bits_source(sinkD_io_d_bits_source),
    .io_d_bits_data(sinkD_io_d_bits_data),
    .io_source(sinkD_io_source),
    .io_way(sinkD_io_way),
    .io_set(sinkD_io_set),
    .io_opcode(sinkD_io_opcode),
    .io_put(sinkD_io_put),
    .io_bs_adr_valid(sinkD_io_bs_adr_valid),
    .io_bs_adr_bits_way(sinkD_io_bs_adr_bits_way),
    .io_bs_adr_bits_set(sinkD_io_bs_adr_bits_set),
    .io_bs_dat_data(sinkD_io_bs_dat_data),
    .io_pb_pop_valid(sinkD_io_pb_pop_valid),
    .io_pb_pop_bits_index(sinkD_io_pb_pop_bits_index),
    .io_pb_beat_data(sinkD_io_pb_beat_data),
    .io_pb_beat_mask(sinkD_io_pb_beat_mask)
  );
  Directory_test directory ( // @[Scheduler.scala 89:25]
    .clock(directory_clock),
    .reset(directory_reset),
    .io_write_ready(directory_io_write_ready),
    .io_write_valid(directory_io_write_valid),
    .io_write_bits_way(directory_io_write_bits_way),
    .io_write_bits_data_tag(directory_io_write_bits_data_tag),
    .io_write_bits_data_valid(directory_io_write_bits_data_valid),
    .io_write_bits_set(directory_io_write_bits_set),
    .io_read_ready(directory_io_read_ready),
    .io_read_valid(directory_io_read_valid),
    .io_read_bits_opcode(directory_io_read_bits_opcode),
    .io_read_bits_source(directory_io_read_bits_source),
    .io_read_bits_tag(directory_io_read_bits_tag),
    .io_read_bits_offset(directory_io_read_bits_offset),
    .io_read_bits_put(directory_io_read_bits_put),
    .io_read_bits_data(directory_io_read_bits_data),
    .io_read_bits_mask(directory_io_read_bits_mask),
    .io_read_bits_set(directory_io_read_bits_set),
    .io_result_valid(directory_io_result_valid),
    .io_result_bits_opcode(directory_io_result_bits_opcode),
    .io_result_bits_source(directory_io_result_bits_source),
    .io_result_bits_tag(directory_io_result_bits_tag),
    .io_result_bits_offset(directory_io_result_bits_offset),
    .io_result_bits_put(directory_io_result_bits_put),
    .io_result_bits_data(directory_io_result_bits_data),
    .io_result_bits_mask(directory_io_result_bits_mask),
    .io_result_bits_set(directory_io_result_bits_set),
    .io_result_bits_hit(directory_io_result_bits_hit),
    .io_result_bits_way(directory_io_result_bits_way)
  );
  BankedStore bankedStore ( // @[Scheduler.scala 91:27]
    .clock(bankedStore_clock),
    .reset(bankedStore_reset),
    .io_sinkD_adr_valid(bankedStore_io_sinkD_adr_valid),
    .io_sinkD_adr_bits_way(bankedStore_io_sinkD_adr_bits_way),
    .io_sinkD_adr_bits_set(bankedStore_io_sinkD_adr_bits_set),
    .io_sinkD_dat_data(bankedStore_io_sinkD_dat_data),
    .io_sourceD_radr_valid(bankedStore_io_sourceD_radr_valid),
    .io_sourceD_radr_bits_way(bankedStore_io_sourceD_radr_bits_way),
    .io_sourceD_radr_bits_set(bankedStore_io_sourceD_radr_bits_set),
    .io_sourceD_radr_bits_mask(bankedStore_io_sourceD_radr_bits_mask),
    .io_sourceD_rdat_data(bankedStore_io_sourceD_rdat_data),
    .io_sourceD_wadr_valid(bankedStore_io_sourceD_wadr_valid),
    .io_sourceD_wadr_bits_way(bankedStore_io_sourceD_wadr_bits_way),
    .io_sourceD_wadr_bits_set(bankedStore_io_sourceD_wadr_bits_set),
    .io_sourceD_wadr_bits_mask(bankedStore_io_sourceD_wadr_bits_mask),
    .io_sourceD_wdat_data(bankedStore_io_sourceD_wdat_data)
  );
  ListBuffer_1 requests ( // @[Scheduler.scala 94:24]
    .clock(requests_clock),
    .reset(requests_reset),
    .io_push_ready(requests_io_push_ready),
    .io_push_valid(requests_io_push_valid),
    .io_push_bits_index(requests_io_push_bits_index),
    .io_push_bits_data(requests_io_push_bits_data),
    .io_valid(requests_io_valid),
    .io_pop_valid(requests_io_pop_valid),
    .io_pop_bits(requests_io_pop_bits),
    .io_data(requests_io_data)
  );
  MSHR_4 mshrs_0 ( // @[Scheduler.scala 96:46]
    .clock(mshrs_0_clock),
    .reset(mshrs_0_reset),
    .io_allocate_valid(mshrs_0_io_allocate_valid),
    .io_allocate_bits_opcode(mshrs_0_io_allocate_bits_opcode),
    .io_allocate_bits_tag(mshrs_0_io_allocate_bits_tag),
    .io_allocate_bits_offset(mshrs_0_io_allocate_bits_offset),
    .io_allocate_bits_put(mshrs_0_io_allocate_bits_put),
    .io_allocate_bits_data(mshrs_0_io_allocate_bits_data),
    .io_allocate_bits_mask(mshrs_0_io_allocate_bits_mask),
    .io_allocate_bits_set(mshrs_0_io_allocate_bits_set),
    .io_allocate_bits_way(mshrs_0_io_allocate_bits_way),
    .io_status_opcode(mshrs_0_io_status_opcode),
    .io_status_tag(mshrs_0_io_status_tag),
    .io_status_put(mshrs_0_io_status_put),
    .io_status_set(mshrs_0_io_status_set),
    .io_status_way(mshrs_0_io_status_way),
    .io_valid(mshrs_0_io_valid),
    .io_schedule_a_ready(mshrs_0_io_schedule_a_ready),
    .io_schedule_a_valid(mshrs_0_io_schedule_a_valid),
    .io_schedule_a_bits_tag(mshrs_0_io_schedule_a_bits_tag),
    .io_schedule_a_bits_offset(mshrs_0_io_schedule_a_bits_offset),
    .io_schedule_a_bits_data(mshrs_0_io_schedule_a_bits_data),
    .io_schedule_a_bits_set(mshrs_0_io_schedule_a_bits_set),
    .io_schedule_d_valid(mshrs_0_io_schedule_d_valid),
    .io_schedule_d_bits_opcode(mshrs_0_io_schedule_d_bits_opcode),
    .io_schedule_d_bits_tag(mshrs_0_io_schedule_d_bits_tag),
    .io_schedule_d_bits_offset(mshrs_0_io_schedule_d_bits_offset),
    .io_schedule_d_bits_put(mshrs_0_io_schedule_d_bits_put),
    .io_schedule_d_bits_data(mshrs_0_io_schedule_d_bits_data),
    .io_schedule_d_bits_mask(mshrs_0_io_schedule_d_bits_mask),
    .io_schedule_d_bits_set(mshrs_0_io_schedule_d_bits_set),
    .io_schedule_d_bits_way(mshrs_0_io_schedule_d_bits_way),
    .io_schedule_dir_ready(mshrs_0_io_schedule_dir_ready),
    .io_schedule_dir_valid(mshrs_0_io_schedule_dir_valid),
    .io_schedule_dir_bits_way(mshrs_0_io_schedule_dir_bits_way),
    .io_schedule_dir_bits_data_tag(mshrs_0_io_schedule_dir_bits_data_tag),
    .io_schedule_dir_bits_set(mshrs_0_io_schedule_dir_bits_set),
    .io_sinkd_valid(mshrs_0_io_sinkd_valid),
    .io_sinkd_bits_data(mshrs_0_io_sinkd_bits_data)
  );
  MSHR_4 mshrs_1 ( // @[Scheduler.scala 96:46]
    .clock(mshrs_1_clock),
    .reset(mshrs_1_reset),
    .io_allocate_valid(mshrs_1_io_allocate_valid),
    .io_allocate_bits_opcode(mshrs_1_io_allocate_bits_opcode),
    .io_allocate_bits_tag(mshrs_1_io_allocate_bits_tag),
    .io_allocate_bits_offset(mshrs_1_io_allocate_bits_offset),
    .io_allocate_bits_put(mshrs_1_io_allocate_bits_put),
    .io_allocate_bits_data(mshrs_1_io_allocate_bits_data),
    .io_allocate_bits_mask(mshrs_1_io_allocate_bits_mask),
    .io_allocate_bits_set(mshrs_1_io_allocate_bits_set),
    .io_allocate_bits_way(mshrs_1_io_allocate_bits_way),
    .io_status_opcode(mshrs_1_io_status_opcode),
    .io_status_tag(mshrs_1_io_status_tag),
    .io_status_put(mshrs_1_io_status_put),
    .io_status_set(mshrs_1_io_status_set),
    .io_status_way(mshrs_1_io_status_way),
    .io_valid(mshrs_1_io_valid),
    .io_schedule_a_ready(mshrs_1_io_schedule_a_ready),
    .io_schedule_a_valid(mshrs_1_io_schedule_a_valid),
    .io_schedule_a_bits_tag(mshrs_1_io_schedule_a_bits_tag),
    .io_schedule_a_bits_offset(mshrs_1_io_schedule_a_bits_offset),
    .io_schedule_a_bits_data(mshrs_1_io_schedule_a_bits_data),
    .io_schedule_a_bits_set(mshrs_1_io_schedule_a_bits_set),
    .io_schedule_d_valid(mshrs_1_io_schedule_d_valid),
    .io_schedule_d_bits_opcode(mshrs_1_io_schedule_d_bits_opcode),
    .io_schedule_d_bits_tag(mshrs_1_io_schedule_d_bits_tag),
    .io_schedule_d_bits_offset(mshrs_1_io_schedule_d_bits_offset),
    .io_schedule_d_bits_put(mshrs_1_io_schedule_d_bits_put),
    .io_schedule_d_bits_data(mshrs_1_io_schedule_d_bits_data),
    .io_schedule_d_bits_mask(mshrs_1_io_schedule_d_bits_mask),
    .io_schedule_d_bits_set(mshrs_1_io_schedule_d_bits_set),
    .io_schedule_d_bits_way(mshrs_1_io_schedule_d_bits_way),
    .io_schedule_dir_ready(mshrs_1_io_schedule_dir_ready),
    .io_schedule_dir_valid(mshrs_1_io_schedule_dir_valid),
    .io_schedule_dir_bits_way(mshrs_1_io_schedule_dir_bits_way),
    .io_schedule_dir_bits_data_tag(mshrs_1_io_schedule_dir_bits_data_tag),
    .io_schedule_dir_bits_set(mshrs_1_io_schedule_dir_bits_set),
    .io_sinkd_valid(mshrs_1_io_sinkd_valid),
    .io_sinkd_bits_data(mshrs_1_io_sinkd_bits_data)
  );
  MSHR_4 mshrs_2 ( // @[Scheduler.scala 96:46]
    .clock(mshrs_2_clock),
    .reset(mshrs_2_reset),
    .io_allocate_valid(mshrs_2_io_allocate_valid),
    .io_allocate_bits_opcode(mshrs_2_io_allocate_bits_opcode),
    .io_allocate_bits_tag(mshrs_2_io_allocate_bits_tag),
    .io_allocate_bits_offset(mshrs_2_io_allocate_bits_offset),
    .io_allocate_bits_put(mshrs_2_io_allocate_bits_put),
    .io_allocate_bits_data(mshrs_2_io_allocate_bits_data),
    .io_allocate_bits_mask(mshrs_2_io_allocate_bits_mask),
    .io_allocate_bits_set(mshrs_2_io_allocate_bits_set),
    .io_allocate_bits_way(mshrs_2_io_allocate_bits_way),
    .io_status_opcode(mshrs_2_io_status_opcode),
    .io_status_tag(mshrs_2_io_status_tag),
    .io_status_put(mshrs_2_io_status_put),
    .io_status_set(mshrs_2_io_status_set),
    .io_status_way(mshrs_2_io_status_way),
    .io_valid(mshrs_2_io_valid),
    .io_schedule_a_ready(mshrs_2_io_schedule_a_ready),
    .io_schedule_a_valid(mshrs_2_io_schedule_a_valid),
    .io_schedule_a_bits_tag(mshrs_2_io_schedule_a_bits_tag),
    .io_schedule_a_bits_offset(mshrs_2_io_schedule_a_bits_offset),
    .io_schedule_a_bits_data(mshrs_2_io_schedule_a_bits_data),
    .io_schedule_a_bits_set(mshrs_2_io_schedule_a_bits_set),
    .io_schedule_d_valid(mshrs_2_io_schedule_d_valid),
    .io_schedule_d_bits_opcode(mshrs_2_io_schedule_d_bits_opcode),
    .io_schedule_d_bits_tag(mshrs_2_io_schedule_d_bits_tag),
    .io_schedule_d_bits_offset(mshrs_2_io_schedule_d_bits_offset),
    .io_schedule_d_bits_put(mshrs_2_io_schedule_d_bits_put),
    .io_schedule_d_bits_data(mshrs_2_io_schedule_d_bits_data),
    .io_schedule_d_bits_mask(mshrs_2_io_schedule_d_bits_mask),
    .io_schedule_d_bits_set(mshrs_2_io_schedule_d_bits_set),
    .io_schedule_d_bits_way(mshrs_2_io_schedule_d_bits_way),
    .io_schedule_dir_ready(mshrs_2_io_schedule_dir_ready),
    .io_schedule_dir_valid(mshrs_2_io_schedule_dir_valid),
    .io_schedule_dir_bits_way(mshrs_2_io_schedule_dir_bits_way),
    .io_schedule_dir_bits_data_tag(mshrs_2_io_schedule_dir_bits_data_tag),
    .io_schedule_dir_bits_set(mshrs_2_io_schedule_dir_bits_set),
    .io_sinkd_valid(mshrs_2_io_sinkd_valid),
    .io_sinkd_bits_data(mshrs_2_io_sinkd_bits_data)
  );
  MSHR_4 mshrs_3 ( // @[Scheduler.scala 96:46]
    .clock(mshrs_3_clock),
    .reset(mshrs_3_reset),
    .io_allocate_valid(mshrs_3_io_allocate_valid),
    .io_allocate_bits_opcode(mshrs_3_io_allocate_bits_opcode),
    .io_allocate_bits_tag(mshrs_3_io_allocate_bits_tag),
    .io_allocate_bits_offset(mshrs_3_io_allocate_bits_offset),
    .io_allocate_bits_put(mshrs_3_io_allocate_bits_put),
    .io_allocate_bits_data(mshrs_3_io_allocate_bits_data),
    .io_allocate_bits_mask(mshrs_3_io_allocate_bits_mask),
    .io_allocate_bits_set(mshrs_3_io_allocate_bits_set),
    .io_allocate_bits_way(mshrs_3_io_allocate_bits_way),
    .io_status_opcode(mshrs_3_io_status_opcode),
    .io_status_tag(mshrs_3_io_status_tag),
    .io_status_put(mshrs_3_io_status_put),
    .io_status_set(mshrs_3_io_status_set),
    .io_status_way(mshrs_3_io_status_way),
    .io_valid(mshrs_3_io_valid),
    .io_schedule_a_ready(mshrs_3_io_schedule_a_ready),
    .io_schedule_a_valid(mshrs_3_io_schedule_a_valid),
    .io_schedule_a_bits_tag(mshrs_3_io_schedule_a_bits_tag),
    .io_schedule_a_bits_offset(mshrs_3_io_schedule_a_bits_offset),
    .io_schedule_a_bits_data(mshrs_3_io_schedule_a_bits_data),
    .io_schedule_a_bits_set(mshrs_3_io_schedule_a_bits_set),
    .io_schedule_d_valid(mshrs_3_io_schedule_d_valid),
    .io_schedule_d_bits_opcode(mshrs_3_io_schedule_d_bits_opcode),
    .io_schedule_d_bits_tag(mshrs_3_io_schedule_d_bits_tag),
    .io_schedule_d_bits_offset(mshrs_3_io_schedule_d_bits_offset),
    .io_schedule_d_bits_put(mshrs_3_io_schedule_d_bits_put),
    .io_schedule_d_bits_data(mshrs_3_io_schedule_d_bits_data),
    .io_schedule_d_bits_mask(mshrs_3_io_schedule_d_bits_mask),
    .io_schedule_d_bits_set(mshrs_3_io_schedule_d_bits_set),
    .io_schedule_d_bits_way(mshrs_3_io_schedule_d_bits_way),
    .io_schedule_dir_ready(mshrs_3_io_schedule_dir_ready),
    .io_schedule_dir_valid(mshrs_3_io_schedule_dir_valid),
    .io_schedule_dir_bits_way(mshrs_3_io_schedule_dir_bits_way),
    .io_schedule_dir_bits_data_tag(mshrs_3_io_schedule_dir_bits_data_tag),
    .io_schedule_dir_bits_set(mshrs_3_io_schedule_dir_bits_set),
    .io_sinkd_valid(mshrs_3_io_sinkd_valid),
    .io_sinkd_bits_data(mshrs_3_io_sinkd_bits_data)
  );
  Queue_106 write_buffer ( // @[Scheduler.scala 140:27]
    .clock(write_buffer_clock),
    .reset(write_buffer_reset),
    .io_enq_ready(write_buffer_io_enq_ready),
    .io_enq_valid(write_buffer_io_enq_valid),
    .io_enq_bits_source(write_buffer_io_enq_bits_source),
    .io_enq_bits_tag(write_buffer_io_enq_bits_tag),
    .io_enq_bits_offset(write_buffer_io_enq_bits_offset),
    .io_enq_bits_data(write_buffer_io_enq_bits_data),
    .io_enq_bits_mask(write_buffer_io_enq_bits_mask),
    .io_enq_bits_set(write_buffer_io_enq_bits_set),
    .io_deq_ready(write_buffer_io_deq_ready),
    .io_deq_valid(write_buffer_io_deq_valid),
    .io_deq_bits_opcode(write_buffer_io_deq_bits_opcode),
    .io_deq_bits_source(write_buffer_io_deq_bits_source),
    .io_deq_bits_tag(write_buffer_io_deq_bits_tag),
    .io_deq_bits_offset(write_buffer_io_deq_bits_offset),
    .io_deq_bits_data(write_buffer_io_deq_bits_data),
    .io_deq_bits_mask(write_buffer_io_deq_bits_mask),
    .io_deq_bits_set(write_buffer_io_deq_bits_set)
  );
  Queue_107 dir_result_buffer ( // @[Scheduler.scala 211:31]
    .clock(dir_result_buffer_clock),
    .reset(dir_result_buffer_reset),
    .io_enq_ready(dir_result_buffer_io_enq_ready),
    .io_enq_valid(dir_result_buffer_io_enq_valid),
    .io_enq_bits_opcode(dir_result_buffer_io_enq_bits_opcode),
    .io_enq_bits_source(dir_result_buffer_io_enq_bits_source),
    .io_enq_bits_tag(dir_result_buffer_io_enq_bits_tag),
    .io_enq_bits_offset(dir_result_buffer_io_enq_bits_offset),
    .io_enq_bits_put(dir_result_buffer_io_enq_bits_put),
    .io_enq_bits_data(dir_result_buffer_io_enq_bits_data),
    .io_enq_bits_mask(dir_result_buffer_io_enq_bits_mask),
    .io_enq_bits_set(dir_result_buffer_io_enq_bits_set),
    .io_enq_bits_hit(dir_result_buffer_io_enq_bits_hit),
    .io_enq_bits_way(dir_result_buffer_io_enq_bits_way),
    .io_deq_ready(dir_result_buffer_io_deq_ready),
    .io_deq_valid(dir_result_buffer_io_deq_valid),
    .io_deq_bits_opcode(dir_result_buffer_io_deq_bits_opcode),
    .io_deq_bits_source(dir_result_buffer_io_deq_bits_source),
    .io_deq_bits_tag(dir_result_buffer_io_deq_bits_tag),
    .io_deq_bits_offset(dir_result_buffer_io_deq_bits_offset),
    .io_deq_bits_put(dir_result_buffer_io_deq_bits_put),
    .io_deq_bits_data(dir_result_buffer_io_deq_bits_data),
    .io_deq_bits_mask(dir_result_buffer_io_deq_bits_mask),
    .io_deq_bits_set(dir_result_buffer_io_deq_bits_set),
    .io_deq_bits_hit(dir_result_buffer_io_deq_bits_hit),
    .io_deq_bits_way(dir_result_buffer_io_deq_bits_way)
  );
  assign io_in_a_ready = sinkA_io_a_ready; // @[Scheduler.scala 79:16]
  assign io_in_d_valid = sourceD_io_d_valid; // @[Scheduler.scala 81:17]
  assign io_in_d_bits_source = sourceD_io_d_bits_source; // @[Scheduler.scala 82:17]
  assign io_in_d_bits_data = sourceD_io_d_bits_data; // @[Scheduler.scala 82:17]
  assign io_in_d_bits_address = sourceD_io_d_bits_address; // @[Scheduler.scala 82:17]
  assign io_out_a_valid = sourceA_io_a_valid; // @[Scheduler.scala 55:18]
  assign io_out_a_bits_opcode = sourceA_io_a_bits_opcode; // @[Scheduler.scala 56:16]
  assign io_out_a_bits_source = sourceA_io_a_bits_source; // @[Scheduler.scala 56:16]
  assign io_out_a_bits_address = sourceA_io_a_bits_address; // @[Scheduler.scala 56:16]
  assign io_out_a_bits_mask = sourceA_io_a_bits_mask; // @[Scheduler.scala 56:16]
  assign io_out_a_bits_data = sourceA_io_a_bits_data; // @[Scheduler.scala 56:16]
  assign io_out_d_ready = sinkD_io_d_ready; // @[Scheduler.scala 67:17]
  assign sourceA_io_req_valid = schedule_a_valid ? schedule_a_valid : write_buffer_io_deq_valid; // @[Scheduler.scala 146:28]
  assign sourceA_io_req_bits_opcode = schedule_a_valid ? schedule_a_bits_opcode : write_buffer_io_deq_bits_opcode; // @[Scheduler.scala 144:27]
  assign sourceA_io_req_bits_source = schedule_a_valid ? schedule_a_bits_source : write_buffer_io_deq_bits_source; // @[Scheduler.scala 144:27]
  assign sourceA_io_req_bits_tag = schedule_a_valid ? schedule_a_bits_tag : write_buffer_io_deq_bits_tag; // @[Scheduler.scala 144:27]
  assign sourceA_io_req_bits_offset = schedule_a_valid ? schedule_a_bits_offset : write_buffer_io_deq_bits_offset; // @[Scheduler.scala 144:27]
  assign sourceA_io_req_bits_data = schedule_a_valid ? schedule_a_bits_data : write_buffer_io_deq_bits_data; // @[Scheduler.scala 144:27]
  assign sourceA_io_req_bits_mask = schedule_a_valid ? schedule_a_bits_mask : write_buffer_io_deq_bits_mask; // @[Scheduler.scala 144:27]
  assign sourceA_io_req_bits_set = schedule_a_valid ? schedule_a_bits_set : write_buffer_io_deq_bits_set; // @[Scheduler.scala 144:27]
  assign sourceA_io_a_ready = io_out_a_ready; // @[Scheduler.scala 57:21]
  assign sourceD_clock = clock;
  assign sourceD_reset = reset;
  assign sourceD_io_req_valid = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_valid : schedule_d_valid; // @[Scheduler.scala 230:28]
  assign sourceD_io_req_bits_opcode = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_opcode :
    schedule_d_bits_opcode; // @[Scheduler.scala 227:34]
  assign sourceD_io_req_bits_source = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_source :
    requests_io_data; // @[Scheduler.scala 231:34]
  assign sourceD_io_req_bits_tag = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_tag :
    schedule_d_bits_tag; // @[Scheduler.scala 224:31]
  assign sourceD_io_req_bits_offset = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_offset :
    schedule_d_bits_offset; // @[Scheduler.scala 226:34]
  assign sourceD_io_req_bits_put = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_put :
    schedule_d_bits_put; // @[Scheduler.scala 228:31]
  assign sourceD_io_req_bits_data = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_data :
    schedule_d_bits_data; // @[Scheduler.scala 220:32]
  assign sourceD_io_req_bits_mask = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_mask :
    schedule_d_bits_mask; // @[Scheduler.scala 225:32]
  assign sourceD_io_req_bits_set = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_set :
    schedule_d_bits_set; // @[Scheduler.scala 223:31]
  assign sourceD_io_req_bits_hit = _dir_result_buffer_io_deq_ready_T & dir_result_buffer_io_deq_bits_hit; // @[Scheduler.scala 222:31]
  assign sourceD_io_req_bits_way = _dir_result_buffer_io_deq_ready_T ? dir_result_buffer_io_deq_bits_way :
    schedule_d_bits_way; // @[Scheduler.scala 219:31]
  assign sourceD_io_req_bits_from_mem = _dir_result_buffer_io_deq_ready_T ? 1'h0 : 1'h1; // @[Scheduler.scala 221:36]
  assign sourceD_io_d_ready = io_in_d_ready; // @[Scheduler.scala 83:21]
  assign sourceD_io_pb_beat_data = sinkA_io_pb_beat_data; // @[Scheduler.scala 63:21]
  assign sourceD_io_pb_beat_mask = sinkA_io_pb_beat_mask; // @[Scheduler.scala 63:21]
  assign sourceD_io_bs_rdat_data = bankedStore_io_sourceD_rdat_data; // @[Scheduler.scala 241:22]
  assign sourceD_io_a_ready = write_buffer_io_enq_ready; // @[Scheduler.scala 147:21]
  assign sinkA_clock = clock;
  assign sinkA_reset = reset;
  assign sinkA_io_req_ready = mshr_free & requests_io_push_ready & (directory_io_read_ready | directory_io_write_ready); // @[Scheduler.scala 206:56]
  assign sinkA_io_a_valid = io_in_a_valid; // @[Scheduler.scala 75:19]
  assign sinkA_io_a_bits_opcode = io_in_a_bits_opcode; // @[Scheduler.scala 74:18]
  assign sinkA_io_a_bits_source = io_in_a_bits_source; // @[Scheduler.scala 74:18]
  assign sinkA_io_a_bits_address = io_in_a_bits_address; // @[Scheduler.scala 74:18]
  assign sinkA_io_a_bits_mask = io_in_a_bits_mask; // @[Scheduler.scala 74:18]
  assign sinkA_io_a_bits_data = io_in_a_bits_data; // @[Scheduler.scala 74:18]
  assign sinkA_io_pb_pop_valid = sourceD_io_pb_pop_valid; // @[Scheduler.scala 62:20]
  assign sinkA_io_pb_pop_bits_index = sourceD_io_pb_pop_bits_index; // @[Scheduler.scala 62:20]
  assign sinkA_io_pb_pop2_valid = sinkD_io_pb_pop_valid; // @[Scheduler.scala 60:19]
  assign sinkA_io_pb_pop2_bits_index = sinkD_io_pb_pop_bits_index; // @[Scheduler.scala 60:19]
  assign sinkD_clock = clock;
  assign sinkD_reset = reset;
  assign sinkD_io_d_valid = io_out_d_valid; // @[Scheduler.scala 66:19]
  assign sinkD_io_d_bits_opcode = io_out_d_bits_opcode; // @[Scheduler.scala 65:18]
  assign sinkD_io_d_bits_source = io_out_d_bits_source; // @[Scheduler.scala 65:18]
  assign sinkD_io_d_bits_data = io_out_d_bits_data; // @[Scheduler.scala 65:18]
  assign sinkD_io_way = 2'h3 == sinkD_io_source[1:0] ? _sinkD_io_way_WIRE_3 : _GEN_2; // @[Scheduler.scala 100:{18,18}]
  assign sinkD_io_set = 2'h3 == sinkD_io_source[1:0] ? mshrs_3_io_status_set : _GEN_6; // @[Scheduler.scala 101:{18,18}]
  assign sinkD_io_opcode = 2'h3 == sinkD_io_source[1:0] ? _sinkD_io_opcode_WIRE_3 : _GEN_10; // @[Scheduler.scala 102:{18,18}]
  assign sinkD_io_put = 2'h3 == sinkD_io_source[1:0] ? _sinkD_io_put_WIRE_3 : _GEN_14; // @[Scheduler.scala 103:{18,18}]
  assign sinkD_io_pb_beat_data = sinkA_io_pb_beat2_data; // @[Scheduler.scala 61:19]
  assign sinkD_io_pb_beat_mask = sinkA_io_pb_beat2_mask; // @[Scheduler.scala 61:19]
  assign directory_clock = clock;
  assign directory_reset = reset;
  assign directory_io_write_valid = mshr_selectOH[0] & mshrs_0_io_schedule_dir_valid | mshr_selectOH[1] &
    mshrs_1_io_schedule_dir_valid | mshr_selectOH[2] & mshrs_2_io_schedule_dir_valid | mshr_selectOH[3] &
    mshrs_3_io_schedule_dir_valid; // @[Mux.scala 27:73]
  assign directory_io_write_bits_way = _schedule_T_30 | _schedule_T_28; // @[Mux.scala 27:73]
  assign directory_io_write_bits_data_tag = _schedule_T_23 | _schedule_T_21; // @[Mux.scala 27:73]
  assign directory_io_write_bits_data_valid = mshr_selectOH[0] | mshr_selectOH[1] | mshr_selectOH[2] | mshr_selectOH[3]; // @[Mux.scala 27:73]
  assign directory_io_write_bits_set = mshr_selectOH[0] & mshrs_0_io_schedule_dir_bits_set | mshr_selectOH[1] &
    mshrs_1_io_schedule_dir_bits_set | mshr_selectOH[2] & mshrs_2_io_schedule_dir_bits_set | mshr_selectOH[3] &
    mshrs_3_io_schedule_dir_bits_set; // @[Mux.scala 27:73]
  assign directory_io_read_valid = sinkA_io_req_valid; // @[Scheduler.scala 151:21 152:17]
  assign directory_io_read_bits_opcode = sinkA_io_req_bits_opcode; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_source = sinkA_io_req_bits_source; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_tag = sinkA_io_req_bits_tag; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_offset = sinkA_io_req_bits_offset; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_put = sinkA_io_req_bits_put; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_data = sinkA_io_req_bits_data; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_mask = sinkA_io_req_bits_mask; // @[Scheduler.scala 151:21 153:16]
  assign directory_io_read_bits_set = sinkA_io_req_bits_set; // @[Scheduler.scala 151:21 153:16]
  assign bankedStore_clock = clock;
  assign bankedStore_reset = reset;
  assign bankedStore_io_sinkD_adr_valid = sinkD_io_bs_adr_valid; // @[Scheduler.scala 235:28]
  assign bankedStore_io_sinkD_adr_bits_way = sinkD_io_bs_adr_bits_way; // @[Scheduler.scala 235:28]
  assign bankedStore_io_sinkD_adr_bits_set = sinkD_io_bs_adr_bits_set; // @[Scheduler.scala 235:28]
  assign bankedStore_io_sinkD_dat_data = sinkD_io_bs_dat_data; // @[Scheduler.scala 237:28]
  assign bankedStore_io_sourceD_radr_valid = sourceD_io_bs_radr_valid; // @[Scheduler.scala 238:31]
  assign bankedStore_io_sourceD_radr_bits_way = sourceD_io_bs_radr_bits_way; // @[Scheduler.scala 238:31]
  assign bankedStore_io_sourceD_radr_bits_set = sourceD_io_bs_radr_bits_set; // @[Scheduler.scala 238:31]
  assign bankedStore_io_sourceD_radr_bits_mask = sourceD_io_bs_radr_bits_mask; // @[Scheduler.scala 238:31]
  assign bankedStore_io_sourceD_wadr_valid = sourceD_io_bs_wadr_valid; // @[Scheduler.scala 239:31]
  assign bankedStore_io_sourceD_wadr_bits_way = sourceD_io_bs_wadr_bits_way; // @[Scheduler.scala 239:31]
  assign bankedStore_io_sourceD_wadr_bits_set = sourceD_io_bs_wadr_bits_set; // @[Scheduler.scala 239:31]
  assign bankedStore_io_sourceD_wadr_bits_mask = sourceD_io_bs_wadr_bits_mask; // @[Scheduler.scala 239:31]
  assign bankedStore_io_sourceD_wdat_data = sourceD_io_bs_wdat_data; // @[Scheduler.scala 240:31]
  assign requests_clock = clock;
  assign requests_reset = reset;
  assign requests_io_push_valid = directory_io_result_valid & _tagMatches_T_3; // @[Scheduler.scala 195:60]
  assign requests_io_push_bits_index = _requests_io_push_bits_index_T_7[1:0]; // @[Scheduler.scala 197:31]
  assign requests_io_push_bits_data = directory_io_result_bits_source; // @[Scheduler.scala 196:31]
  assign requests_io_pop_valid = _requests_io_pop_valid_T[0] & schedule_d_valid & sourceD_io_req_ready; // @[Scheduler.scala 202:76]
  assign requests_io_pop_bits = {_mshr_select_T,_mshr_select_T_1[1]}; // @[Cat.scala 31:58]
  assign mshrs_0_clock = clock;
  assign mshrs_0_reset = reset;
  assign mshrs_0_io_allocate_valid = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3; // @[Scheduler.scala 189:51]
  assign mshrs_0_io_allocate_bits_opcode = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_opcode : 3'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_tag = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_tag : 26'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_offset = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_offset : 5'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_put = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_put : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_data = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_data : 256'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_mask = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_mask : 8'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_set = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 &
    directory_io_result_bits_set; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_allocate_bits_way = directory_io_result_valid & alloc & mshr_insertOH[0] & _tagMatches_T_3 ?
    directory_io_result_bits_way : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_0_io_valid = requests_io_valid[0]; // @[Scheduler.scala 135:41]
  assign mshrs_0_io_schedule_a_ready = sourceA_io_req_ready & mshr_select == 2'h0; // @[Scheduler.scala 132:51]
  assign mshrs_0_io_schedule_dir_ready = directory_io_write_ready & _mshrs_0_io_schedule_a_ready_T; // @[Scheduler.scala 134:55]
  assign mshrs_0_io_sinkd_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h0 & sinkD_io_resp_bits_opcode
     == 3'h1; // @[Scheduler.scala 130:90]
  assign mshrs_0_io_sinkd_bits_data = sinkD_io_resp_bits_data; // @[Scheduler.scala 131:22]
  assign mshrs_1_clock = clock;
  assign mshrs_1_reset = reset;
  assign mshrs_1_io_allocate_valid = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3; // @[Scheduler.scala 189:51]
  assign mshrs_1_io_allocate_bits_opcode = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_opcode : 3'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_tag = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_tag : 26'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_offset = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_offset : 5'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_put = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_put : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_data = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_data : 256'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_mask = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_mask : 8'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_set = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 &
    directory_io_result_bits_set; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_allocate_bits_way = directory_io_result_valid & alloc & mshr_insertOH[1] & _tagMatches_T_3 ?
    directory_io_result_bits_way : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_1_io_valid = requests_io_valid[1]; // @[Scheduler.scala 135:41]
  assign mshrs_1_io_schedule_a_ready = sourceA_io_req_ready & mshr_select == 2'h1; // @[Scheduler.scala 132:51]
  assign mshrs_1_io_schedule_dir_ready = directory_io_write_ready & _mshrs_1_io_schedule_a_ready_T; // @[Scheduler.scala 134:55]
  assign mshrs_1_io_sinkd_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h1 & sinkD_io_resp_bits_opcode
     == 3'h1; // @[Scheduler.scala 130:90]
  assign mshrs_1_io_sinkd_bits_data = sinkD_io_resp_bits_data; // @[Scheduler.scala 131:22]
  assign mshrs_2_clock = clock;
  assign mshrs_2_reset = reset;
  assign mshrs_2_io_allocate_valid = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3; // @[Scheduler.scala 189:51]
  assign mshrs_2_io_allocate_bits_opcode = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_opcode : 3'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_tag = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_tag : 26'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_offset = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_offset : 5'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_put = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_put : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_data = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_data : 256'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_mask = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_mask : 8'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_set = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 &
    directory_io_result_bits_set; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_allocate_bits_way = directory_io_result_valid & alloc & mshr_insertOH[2] & _tagMatches_T_3 ?
    directory_io_result_bits_way : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_2_io_valid = requests_io_valid[2]; // @[Scheduler.scala 135:41]
  assign mshrs_2_io_schedule_a_ready = sourceA_io_req_ready & mshr_select == 2'h2; // @[Scheduler.scala 132:51]
  assign mshrs_2_io_schedule_dir_ready = directory_io_write_ready & _mshrs_2_io_schedule_a_ready_T; // @[Scheduler.scala 134:55]
  assign mshrs_2_io_sinkd_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h2 & sinkD_io_resp_bits_opcode
     == 3'h1; // @[Scheduler.scala 130:90]
  assign mshrs_2_io_sinkd_bits_data = sinkD_io_resp_bits_data; // @[Scheduler.scala 131:22]
  assign mshrs_3_clock = clock;
  assign mshrs_3_reset = reset;
  assign mshrs_3_io_allocate_valid = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3; // @[Scheduler.scala 189:51]
  assign mshrs_3_io_allocate_bits_opcode = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_opcode : 3'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_tag = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_tag : 26'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_offset = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_offset : 5'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_put = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_put : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_data = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_data : 256'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_mask = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_mask : 8'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_set = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 &
    directory_io_result_bits_set; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_allocate_bits_way = directory_io_result_valid & alloc & mshr_insertOH[3] & _tagMatches_T_3 ?
    directory_io_result_bits_way : 2'h0; // @[Scheduler.scala 188:23 189:84 191:26]
  assign mshrs_3_io_valid = requests_io_valid[3]; // @[Scheduler.scala 135:41]
  assign mshrs_3_io_schedule_a_ready = sourceA_io_req_ready & mshr_select == 2'h3; // @[Scheduler.scala 132:51]
  assign mshrs_3_io_schedule_dir_ready = directory_io_write_ready & _mshrs_3_io_schedule_a_ready_T; // @[Scheduler.scala 134:55]
  assign mshrs_3_io_sinkd_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h3 & sinkD_io_resp_bits_opcode
     == 3'h1; // @[Scheduler.scala 130:90]
  assign mshrs_3_io_sinkd_bits_data = sinkD_io_resp_bits_data; // @[Scheduler.scala 131:22]
  assign write_buffer_clock = clock;
  assign write_buffer_reset = reset;
  assign write_buffer_io_enq_valid = sourceD_io_a_valid; // @[Scheduler.scala 141:28]
  assign write_buffer_io_enq_bits_source = sourceD_io_a_bits_source; // @[Scheduler.scala 142:27]
  assign write_buffer_io_enq_bits_tag = sourceD_io_a_bits_tag; // @[Scheduler.scala 142:27]
  assign write_buffer_io_enq_bits_offset = sourceD_io_a_bits_offset; // @[Scheduler.scala 142:27]
  assign write_buffer_io_enq_bits_data = sourceD_io_a_bits_data; // @[Scheduler.scala 142:27]
  assign write_buffer_io_enq_bits_mask = sourceD_io_a_bits_mask; // @[Scheduler.scala 142:27]
  assign write_buffer_io_enq_bits_set = sourceD_io_a_bits_set; // @[Scheduler.scala 142:27]
  assign write_buffer_io_deq_ready = sourceA_io_req_ready & ~schedule_a_valid; // @[Scheduler.scala 143:51]
  assign dir_result_buffer_clock = clock;
  assign dir_result_buffer_reset = reset;
  assign dir_result_buffer_io_enq_valid = directory_io_result_valid & directory_io_result_bits_hit; // @[Scheduler.scala 213:62]
  assign dir_result_buffer_io_enq_bits_opcode = directory_io_result_bits_opcode; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_source = directory_io_result_bits_source; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_offset = directory_io_result_bits_offset; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_put = directory_io_result_bits_put; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_data = directory_io_result_bits_data; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_mask = directory_io_result_bits_mask; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_set = directory_io_result_bits_set; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_enq_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 214:32]
  assign dir_result_buffer_io_deq_ready = ~schedule_d_valid; // @[Scheduler.scala 215:36]
  always @(posedge clock) begin
    if (reset) begin // @[Scheduler.scala 113:29]
      robin_filter <= 4'h0; // @[Scheduler.scala 113:29]
    end else if (|mshr_request) begin // @[Scheduler.scala 124:29]
      robin_filter <= _robin_filter_T_5; // @[Scheduler.scala 124:44]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  robin_filter = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_32(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [2:0]   io_in_0_bits_opcode,
  input  [3:0]   io_in_0_bits_source,
  input  [31:0]  io_in_0_bits_address,
  input  [31:0]  io_in_0_bits_mask,
  input  [255:0] io_in_0_bits_data,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [2:0]   io_in_1_bits_opcode,
  input  [3:0]   io_in_1_bits_source,
  input  [31:0]  io_in_1_bits_address,
  input  [31:0]  io_in_1_bits_mask,
  input  [255:0] io_in_1_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_opcode,
  output [3:0]   io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [31:0]  io_out_bits_mask,
  output [255:0] io_out_bits_data
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 46:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 149:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 149:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_opcode = io_in_0_valid ? io_in_0_bits_opcode : io_in_1_bits_opcode; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_source = io_in_0_valid ? io_in_0_bits_source : io_in_1_bits_source; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_address = io_in_0_valid ? io_in_0_bits_address : io_in_1_bits_address; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_mask = io_in_0_valid ? io_in_0_bits_mask : io_in_1_bits_mask; // @[Arbiter.scala 139:15 141:26 143:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 139:15 141:26 143:19]
endmodule
module SM2L2Arbiter(
  output         io_memReqVecIn_0_ready,
  input          io_memReqVecIn_0_valid,
  input  [2:0]   io_memReqVecIn_0_bits_a_opcode,
  input  [31:0]  io_memReqVecIn_0_bits_a_addr,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_0,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_1,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_2,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_3,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_4,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_5,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_6,
  input  [31:0]  io_memReqVecIn_0_bits_a_data_7,
  input          io_memReqVecIn_0_bits_a_mask_0,
  input          io_memReqVecIn_0_bits_a_mask_1,
  input          io_memReqVecIn_0_bits_a_mask_2,
  input          io_memReqVecIn_0_bits_a_mask_3,
  input          io_memReqVecIn_0_bits_a_mask_4,
  input          io_memReqVecIn_0_bits_a_mask_5,
  input          io_memReqVecIn_0_bits_a_mask_6,
  input          io_memReqVecIn_0_bits_a_mask_7,
  input  [2:0]   io_memReqVecIn_0_bits_a_source,
  output         io_memReqVecIn_1_ready,
  input          io_memReqVecIn_1_valid,
  input  [2:0]   io_memReqVecIn_1_bits_a_opcode,
  input  [31:0]  io_memReqVecIn_1_bits_a_addr,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_0,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_1,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_2,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_3,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_4,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_5,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_6,
  input  [31:0]  io_memReqVecIn_1_bits_a_data_7,
  input          io_memReqVecIn_1_bits_a_mask_0,
  input          io_memReqVecIn_1_bits_a_mask_1,
  input          io_memReqVecIn_1_bits_a_mask_2,
  input          io_memReqVecIn_1_bits_a_mask_3,
  input          io_memReqVecIn_1_bits_a_mask_4,
  input          io_memReqVecIn_1_bits_a_mask_5,
  input          io_memReqVecIn_1_bits_a_mask_6,
  input          io_memReqVecIn_1_bits_a_mask_7,
  input  [2:0]   io_memReqVecIn_1_bits_a_source,
  input          io_memReqOut_ready,
  output         io_memReqOut_valid,
  output [2:0]   io_memReqOut_bits_opcode,
  output [3:0]   io_memReqOut_bits_source,
  output [31:0]  io_memReqOut_bits_address,
  output [31:0]  io_memReqOut_bits_mask,
  output [255:0] io_memReqOut_bits_data,
  output         io_memRspIn_ready,
  input          io_memRspIn_valid,
  input  [3:0]   io_memRspIn_bits_source,
  input  [255:0] io_memRspIn_bits_data,
  input  [31:0]  io_memRspIn_bits_address,
  input          io_memRspVecOut_0_ready,
  output         io_memRspVecOut_0_valid,
  output [31:0]  io_memRspVecOut_0_bits_d_addr,
  output [31:0]  io_memRspVecOut_0_bits_d_data_0,
  output [31:0]  io_memRspVecOut_0_bits_d_data_1,
  output [31:0]  io_memRspVecOut_0_bits_d_data_2,
  output [31:0]  io_memRspVecOut_0_bits_d_data_3,
  output [31:0]  io_memRspVecOut_0_bits_d_data_4,
  output [31:0]  io_memRspVecOut_0_bits_d_data_5,
  output [31:0]  io_memRspVecOut_0_bits_d_data_6,
  output [31:0]  io_memRspVecOut_0_bits_d_data_7,
  output [2:0]   io_memRspVecOut_0_bits_d_source,
  input          io_memRspVecOut_1_ready,
  output         io_memRspVecOut_1_valid,
  output [31:0]  io_memRspVecOut_1_bits_d_addr,
  output [31:0]  io_memRspVecOut_1_bits_d_data_0,
  output [31:0]  io_memRspVecOut_1_bits_d_data_1,
  output [31:0]  io_memRspVecOut_1_bits_d_data_2,
  output [31:0]  io_memRspVecOut_1_bits_d_data_3,
  output [31:0]  io_memRspVecOut_1_bits_d_data_4,
  output [31:0]  io_memRspVecOut_1_bits_d_data_5,
  output [31:0]  io_memRspVecOut_1_bits_d_data_6,
  output [31:0]  io_memRspVecOut_1_bits_d_data_7,
  output [2:0]   io_memRspVecOut_1_bits_d_source
);
  wire  memReqArb_io_in_0_ready; // @[GPGPU_top.scala 252:25]
  wire  memReqArb_io_in_0_valid; // @[GPGPU_top.scala 252:25]
  wire [2:0] memReqArb_io_in_0_bits_opcode; // @[GPGPU_top.scala 252:25]
  wire [3:0] memReqArb_io_in_0_bits_source; // @[GPGPU_top.scala 252:25]
  wire [31:0] memReqArb_io_in_0_bits_address; // @[GPGPU_top.scala 252:25]
  wire [31:0] memReqArb_io_in_0_bits_mask; // @[GPGPU_top.scala 252:25]
  wire [255:0] memReqArb_io_in_0_bits_data; // @[GPGPU_top.scala 252:25]
  wire  memReqArb_io_in_1_ready; // @[GPGPU_top.scala 252:25]
  wire  memReqArb_io_in_1_valid; // @[GPGPU_top.scala 252:25]
  wire [2:0] memReqArb_io_in_1_bits_opcode; // @[GPGPU_top.scala 252:25]
  wire [3:0] memReqArb_io_in_1_bits_source; // @[GPGPU_top.scala 252:25]
  wire [31:0] memReqArb_io_in_1_bits_address; // @[GPGPU_top.scala 252:25]
  wire [31:0] memReqArb_io_in_1_bits_mask; // @[GPGPU_top.scala 252:25]
  wire [255:0] memReqArb_io_in_1_bits_data; // @[GPGPU_top.scala 252:25]
  wire  memReqArb_io_out_ready; // @[GPGPU_top.scala 252:25]
  wire  memReqArb_io_out_valid; // @[GPGPU_top.scala 252:25]
  wire [2:0] memReqArb_io_out_bits_opcode; // @[GPGPU_top.scala 252:25]
  wire [3:0] memReqArb_io_out_bits_source; // @[GPGPU_top.scala 252:25]
  wire [31:0] memReqArb_io_out_bits_address; // @[GPGPU_top.scala 252:25]
  wire [31:0] memReqArb_io_out_bits_mask; // @[GPGPU_top.scala 252:25]
  wire [255:0] memReqArb_io_out_bits_data; // @[GPGPU_top.scala 252:25]
  wire [7:0] _memReqArb_io_in_0_bits_mask_T = {io_memReqVecIn_0_bits_a_mask_7,io_memReqVecIn_0_bits_a_mask_6,
    io_memReqVecIn_0_bits_a_mask_5,io_memReqVecIn_0_bits_a_mask_4,io_memReqVecIn_0_bits_a_mask_3,
    io_memReqVecIn_0_bits_a_mask_2,io_memReqVecIn_0_bits_a_mask_1,io_memReqVecIn_0_bits_a_mask_0}; // @[GPGPU_top.scala 258:69]
  wire [127:0] memReqArb_io_in_0_bits_data_lo = {io_memReqVecIn_0_bits_a_data_3,io_memReqVecIn_0_bits_a_data_2,
    io_memReqVecIn_0_bits_a_data_1,io_memReqVecIn_0_bits_a_data_0}; // @[GPGPU_top.scala 259:67]
  wire [127:0] memReqArb_io_in_0_bits_data_hi = {io_memReqVecIn_0_bits_a_data_7,io_memReqVecIn_0_bits_a_data_6,
    io_memReqVecIn_0_bits_a_data_5,io_memReqVecIn_0_bits_a_data_4}; // @[GPGPU_top.scala 259:67]
  wire [7:0] _memReqArb_io_in_1_bits_mask_T = {io_memReqVecIn_1_bits_a_mask_7,io_memReqVecIn_1_bits_a_mask_6,
    io_memReqVecIn_1_bits_a_mask_5,io_memReqVecIn_1_bits_a_mask_4,io_memReqVecIn_1_bits_a_mask_3,
    io_memReqVecIn_1_bits_a_mask_2,io_memReqVecIn_1_bits_a_mask_1,io_memReqVecIn_1_bits_a_mask_0}; // @[GPGPU_top.scala 258:69]
  wire [127:0] memReqArb_io_in_1_bits_data_lo = {io_memReqVecIn_1_bits_a_data_3,io_memReqVecIn_1_bits_a_data_2,
    io_memReqVecIn_1_bits_a_data_1,io_memReqVecIn_1_bits_a_data_0}; // @[GPGPU_top.scala 259:67]
  wire [127:0] memReqArb_io_in_1_bits_data_hi = {io_memReqVecIn_1_bits_a_data_7,io_memReqVecIn_1_bits_a_data_6,
    io_memReqVecIn_1_bits_a_data_5,io_memReqVecIn_1_bits_a_data_4}; // @[GPGPU_top.scala 259:67]
  wire [1:0] _io_memRspIn_ready_T_1 = 2'h1 << io_memRspIn_bits_source[3]; // @[OneHot.scala 57:35]
  wire [1:0] _io_memRspIn_ready_T_2 = {io_memRspVecOut_0_ready,io_memRspVecOut_1_ready}; // @[Cat.scala 31:58]
  wire [1:0] _io_memRspIn_ready_T_5 = {_io_memRspIn_ready_T_2[0],_io_memRspIn_ready_T_2[1]}; // @[Cat.scala 31:58]
  wire [1:0] _io_memRspIn_ready_T_6 = _io_memRspIn_ready_T_1 & _io_memRspIn_ready_T_5; // @[Mux.scala 30:47]
  Arbiter_32 memReqArb ( // @[GPGPU_top.scala 252:25]
    .io_in_0_ready(memReqArb_io_in_0_ready),
    .io_in_0_valid(memReqArb_io_in_0_valid),
    .io_in_0_bits_opcode(memReqArb_io_in_0_bits_opcode),
    .io_in_0_bits_source(memReqArb_io_in_0_bits_source),
    .io_in_0_bits_address(memReqArb_io_in_0_bits_address),
    .io_in_0_bits_mask(memReqArb_io_in_0_bits_mask),
    .io_in_0_bits_data(memReqArb_io_in_0_bits_data),
    .io_in_1_ready(memReqArb_io_in_1_ready),
    .io_in_1_valid(memReqArb_io_in_1_valid),
    .io_in_1_bits_opcode(memReqArb_io_in_1_bits_opcode),
    .io_in_1_bits_source(memReqArb_io_in_1_bits_source),
    .io_in_1_bits_address(memReqArb_io_in_1_bits_address),
    .io_in_1_bits_mask(memReqArb_io_in_1_bits_mask),
    .io_in_1_bits_data(memReqArb_io_in_1_bits_data),
    .io_out_ready(memReqArb_io_out_ready),
    .io_out_valid(memReqArb_io_out_valid),
    .io_out_bits_opcode(memReqArb_io_out_bits_opcode),
    .io_out_bits_source(memReqArb_io_out_bits_source),
    .io_out_bits_address(memReqArb_io_out_bits_address),
    .io_out_bits_mask(memReqArb_io_out_bits_mask),
    .io_out_bits_data(memReqArb_io_out_bits_data)
  );
  assign io_memReqVecIn_0_ready = memReqArb_io_in_0_ready; // @[GPGPU_top.scala 262:28]
  assign io_memReqVecIn_1_ready = memReqArb_io_in_1_ready; // @[GPGPU_top.scala 262:28]
  assign io_memReqOut_valid = memReqArb_io_out_valid; // @[GPGPU_top.scala 264:16]
  assign io_memReqOut_bits_opcode = memReqArb_io_out_bits_opcode; // @[GPGPU_top.scala 264:16]
  assign io_memReqOut_bits_source = memReqArb_io_out_bits_source; // @[GPGPU_top.scala 264:16]
  assign io_memReqOut_bits_address = memReqArb_io_out_bits_address; // @[GPGPU_top.scala 264:16]
  assign io_memReqOut_bits_mask = memReqArb_io_out_bits_mask; // @[GPGPU_top.scala 264:16]
  assign io_memReqOut_bits_data = memReqArb_io_out_bits_data; // @[GPGPU_top.scala 264:16]
  assign io_memRspIn_ready = |_io_memRspIn_ready_T_6; // @[Mux.scala 30:53]
  assign io_memRspVecOut_0_valid = ~io_memRspIn_bits_source[3] & io_memRspIn_valid; // @[GPGPU_top.scala 273:112]
  assign io_memRspVecOut_0_bits_d_addr = io_memRspIn_bits_address; // @[GPGPU_top.scala 271:35]
  assign io_memRspVecOut_0_bits_d_data_0 = io_memRspIn_bits_data[31:0]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_1 = io_memRspIn_bits_data[63:32]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_2 = io_memRspIn_bits_data[95:64]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_3 = io_memRspIn_bits_data[127:96]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_4 = io_memRspIn_bits_data[159:128]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_5 = io_memRspIn_bits_data[191:160]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_6 = io_memRspIn_bits_data[223:192]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_data_7 = io_memRspIn_bits_data[255:224]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_0_bits_d_source = io_memRspIn_bits_source[2:0]; // @[GPGPU_top.scala 270:37]
  assign io_memRspVecOut_1_valid = io_memRspIn_bits_source[3] & io_memRspIn_valid; // @[GPGPU_top.scala 273:112]
  assign io_memRspVecOut_1_bits_d_addr = io_memRspIn_bits_address; // @[GPGPU_top.scala 271:35]
  assign io_memRspVecOut_1_bits_d_data_0 = io_memRspIn_bits_data[31:0]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_1 = io_memRspIn_bits_data[63:32]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_2 = io_memRspIn_bits_data[95:64]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_3 = io_memRspIn_bits_data[127:96]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_4 = io_memRspIn_bits_data[159:128]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_5 = io_memRspIn_bits_data[191:160]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_6 = io_memRspIn_bits_data[223:192]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_data_7 = io_memRspIn_bits_data[255:224]; // @[GPGPU_top.scala 269:67]
  assign io_memRspVecOut_1_bits_d_source = io_memRspIn_bits_source[2:0]; // @[GPGPU_top.scala 270:37]
  assign memReqArb_io_in_0_valid = io_memReqVecIn_0_valid; // @[GPGPU_top.scala 261:30]
  assign memReqArb_io_in_0_bits_opcode = io_memReqVecIn_0_bits_a_opcode; // @[GPGPU_top.scala 255:36]
  assign memReqArb_io_in_0_bits_source = {1'h0,io_memReqVecIn_0_bits_a_source}; // @[Cat.scala 31:58]
  assign memReqArb_io_in_0_bits_address = io_memReqVecIn_0_bits_a_addr; // @[GPGPU_top.scala 257:37]
  assign memReqArb_io_in_0_bits_mask = {{24'd0}, _memReqArb_io_in_0_bits_mask_T}; // @[GPGPU_top.scala 258:34]
  assign memReqArb_io_in_0_bits_data = {memReqArb_io_in_0_bits_data_hi,memReqArb_io_in_0_bits_data_lo}; // @[GPGPU_top.scala 259:67]
  assign memReqArb_io_in_1_valid = io_memReqVecIn_1_valid; // @[GPGPU_top.scala 261:30]
  assign memReqArb_io_in_1_bits_opcode = io_memReqVecIn_1_bits_a_opcode; // @[GPGPU_top.scala 255:36]
  assign memReqArb_io_in_1_bits_source = {1'h1,io_memReqVecIn_1_bits_a_source}; // @[Cat.scala 31:58]
  assign memReqArb_io_in_1_bits_address = io_memReqVecIn_1_bits_a_addr; // @[GPGPU_top.scala 257:37]
  assign memReqArb_io_in_1_bits_mask = {{24'd0}, _memReqArb_io_in_1_bits_mask_T}; // @[GPGPU_top.scala 258:34]
  assign memReqArb_io_in_1_bits_data = {memReqArb_io_in_1_bits_data_hi,memReqArb_io_in_1_bits_data_lo}; // @[GPGPU_top.scala 259:67]
  assign memReqArb_io_out_ready = io_memReqOut_ready; // @[GPGPU_top.scala 264:16]
endmodule
module GPGPU_top(
  input          clock,
  input          reset,
  output         io_host_req_ready,
  input          io_host_req_valid,
  input  [4:0]   io_host_req_bits_host_wg_id,
  input  [2:0]   io_host_req_bits_host_num_wf,
  input  [9:0]   io_host_req_bits_host_wf_size,
  input  [31:0]  io_host_req_bits_host_start_pc,
  input  [12:0]  io_host_req_bits_host_vgpr_size_total,
  input  [12:0]  io_host_req_bits_host_sgpr_size_total,
  input  [12:0]  io_host_req_bits_host_lds_size_total,
  input  [10:0]  io_host_req_bits_host_gds_size_total,
  input  [12:0]  io_host_req_bits_host_vgpr_size_per_wf,
  input  [12:0]  io_host_req_bits_host_sgpr_size_per_wf,
  input          io_host_rsp_ready,
  output         io_host_rsp_valid,
  output [4:0]   io_host_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id,
  input          io_out_a_ready,
  output         io_out_a_valid,
  output [2:0]   io_out_a_bits_opcode,
  output [3:0]   io_out_a_bits_source,
  output [31:0]  io_out_a_bits_address,
  output [31:0]  io_out_a_bits_mask,
  output [255:0] io_out_a_bits_data,
  output         io_out_d_ready,
  input          io_out_d_valid,
  input  [2:0]   io_out_d_bits_opcode,
  input  [3:0]   io_out_d_bits_source,
  input  [255:0] io_out_d_bits_data
);
  wire  cta_clock; // @[GPGPU_top.scala 116:19]
  wire  cta_reset; // @[GPGPU_top.scala 116:19]
  wire  cta_io_host2CTA_ready; // @[GPGPU_top.scala 116:19]
  wire  cta_io_host2CTA_valid; // @[GPGPU_top.scala 116:19]
  wire [4:0] cta_io_host2CTA_bits_host_wg_id; // @[GPGPU_top.scala 116:19]
  wire [2:0] cta_io_host2CTA_bits_host_num_wf; // @[GPGPU_top.scala 116:19]
  wire [9:0] cta_io_host2CTA_bits_host_wf_size; // @[GPGPU_top.scala 116:19]
  wire [31:0] cta_io_host2CTA_bits_host_start_pc; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_host2CTA_bits_host_vgpr_size_total; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_host2CTA_bits_host_sgpr_size_total; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_host2CTA_bits_host_lds_size_total; // @[GPGPU_top.scala 116:19]
  wire [10:0] cta_io_host2CTA_bits_host_gds_size_total; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_host2CTA_bits_host_vgpr_size_per_wf; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_host2CTA_bits_host_sgpr_size_per_wf; // @[GPGPU_top.scala 116:19]
  wire  cta_io_CTA2host_ready; // @[GPGPU_top.scala 116:19]
  wire  cta_io_CTA2host_valid; // @[GPGPU_top.scala 116:19]
  wire [4:0] cta_io_CTA2host_bits_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 116:19]
  wire  cta_io_CTA2warp_0_ready; // @[GPGPU_top.scala 116:19]
  wire  cta_io_CTA2warp_0_valid; // @[GPGPU_top.scala 116:19]
  wire [2:0] cta_io_CTA2warp_0_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 116:19]
  wire [9:0] cta_io_CTA2warp_0_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_CTA2warp_0_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_CTA2warp_0_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 116:19]
  wire [4:0] cta_io_CTA2warp_0_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_CTA2warp_0_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 116:19]
  wire [31:0] cta_io_CTA2warp_0_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 116:19]
  wire  cta_io_CTA2warp_1_ready; // @[GPGPU_top.scala 116:19]
  wire  cta_io_CTA2warp_1_valid; // @[GPGPU_top.scala 116:19]
  wire [2:0] cta_io_CTA2warp_1_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 116:19]
  wire [9:0] cta_io_CTA2warp_1_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_CTA2warp_1_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_CTA2warp_1_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 116:19]
  wire [4:0] cta_io_CTA2warp_1_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 116:19]
  wire [12:0] cta_io_CTA2warp_1_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 116:19]
  wire [31:0] cta_io_CTA2warp_1_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 116:19]
  wire  cta_io_warp2CTA_0_valid; // @[GPGPU_top.scala 116:19]
  wire [4:0] cta_io_warp2CTA_0_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 116:19]
  wire  cta_io_warp2CTA_1_valid; // @[GPGPU_top.scala 116:19]
  wire [4:0] cta_io_warp2CTA_1_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 116:19]
  wire  SM_wrapper_clock; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_reset; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_CTAreq_ready; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_CTAreq_valid; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 117:47]
  wire [9:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 117:47]
  wire [12:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 117:47]
  wire [12:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 117:47]
  wire [4:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 117:47]
  wire [12:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_CTAreq_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_CTArsp_valid; // @[GPGPU_top.scala 117:47]
  wire [4:0] SM_wrapper_io_CTArsp_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memRsp_ready; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memRsp_valid; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_addr; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_0; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_1; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_2; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_3; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_4; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_5; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_6; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memRsp_bits_d_data_7; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_io_memRsp_bits_d_source; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_ready; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_valid; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_io_memReq_bits_a_opcode; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_addr; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_0; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_1; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_2; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_3; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_4; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_5; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_6; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_io_memReq_bits_a_data_7; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_0; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_1; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_2; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_3; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_4; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_5; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_6; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_io_memReq_bits_a_mask_7; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_io_memReq_bits_a_source; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_clock; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_reset; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_CTAreq_ready; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_CTAreq_valid; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 117:47]
  wire [9:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 117:47]
  wire [12:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 117:47]
  wire [12:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 117:47]
  wire [4:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 117:47]
  wire [12:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_CTAreq_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_CTArsp_valid; // @[GPGPU_top.scala 117:47]
  wire [4:0] SM_wrapper_1_io_CTArsp_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memRsp_ready; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memRsp_valid; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_addr; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_0; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_1; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_2; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_3; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_4; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_5; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_6; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memRsp_bits_d_data_7; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_1_io_memRsp_bits_d_source; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_ready; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_valid; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_1_io_memReq_bits_a_opcode; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_addr; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_0; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_1; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_2; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_3; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_4; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_5; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_6; // @[GPGPU_top.scala 117:47]
  wire [31:0] SM_wrapper_1_io_memReq_bits_a_data_7; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_0; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_1; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_2; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_3; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_4; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_5; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_6; // @[GPGPU_top.scala 117:47]
  wire  SM_wrapper_1_io_memReq_bits_a_mask_7; // @[GPGPU_top.scala 117:47]
  wire [2:0] SM_wrapper_1_io_memReq_bits_a_source; // @[GPGPU_top.scala 117:47]
  wire  l2cache_clock; // @[GPGPU_top.scala 118:21]
  wire  l2cache_reset; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_in_a_ready; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_in_a_valid; // @[GPGPU_top.scala 118:21]
  wire [2:0] l2cache_io_in_a_bits_opcode; // @[GPGPU_top.scala 118:21]
  wire [3:0] l2cache_io_in_a_bits_source; // @[GPGPU_top.scala 118:21]
  wire [31:0] l2cache_io_in_a_bits_address; // @[GPGPU_top.scala 118:21]
  wire [31:0] l2cache_io_in_a_bits_mask; // @[GPGPU_top.scala 118:21]
  wire [255:0] l2cache_io_in_a_bits_data; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_in_d_ready; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_in_d_valid; // @[GPGPU_top.scala 118:21]
  wire [3:0] l2cache_io_in_d_bits_source; // @[GPGPU_top.scala 118:21]
  wire [255:0] l2cache_io_in_d_bits_data; // @[GPGPU_top.scala 118:21]
  wire [31:0] l2cache_io_in_d_bits_address; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_out_a_ready; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_out_a_valid; // @[GPGPU_top.scala 118:21]
  wire [2:0] l2cache_io_out_a_bits_opcode; // @[GPGPU_top.scala 118:21]
  wire [3:0] l2cache_io_out_a_bits_source; // @[GPGPU_top.scala 118:21]
  wire [31:0] l2cache_io_out_a_bits_address; // @[GPGPU_top.scala 118:21]
  wire [31:0] l2cache_io_out_a_bits_mask; // @[GPGPU_top.scala 118:21]
  wire [255:0] l2cache_io_out_a_bits_data; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_out_d_ready; // @[GPGPU_top.scala 118:21]
  wire  l2cache_io_out_d_valid; // @[GPGPU_top.scala 118:21]
  wire [2:0] l2cache_io_out_d_bits_opcode; // @[GPGPU_top.scala 118:21]
  wire [3:0] l2cache_io_out_d_bits_source; // @[GPGPU_top.scala 118:21]
  wire [255:0] l2cache_io_out_d_bits_data; // @[GPGPU_top.scala 118:21]
  wire  sm2L2Arb_io_memReqVecIn_0_ready; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_valid; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memReqVecIn_0_bits_a_opcode; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_addr; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_0; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_1; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_2; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_3; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_4; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_5; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_6; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_0_bits_a_data_7; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_0; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_1; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_2; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_3; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_4; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_5; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_6; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_0_bits_a_mask_7; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memReqVecIn_0_bits_a_source; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_ready; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_valid; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memReqVecIn_1_bits_a_opcode; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_addr; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_0; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_1; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_2; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_3; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_4; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_5; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_6; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqVecIn_1_bits_a_data_7; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_0; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_1; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_2; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_3; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_4; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_5; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_6; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqVecIn_1_bits_a_mask_7; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memReqVecIn_1_bits_a_source; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqOut_ready; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memReqOut_valid; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memReqOut_bits_opcode; // @[GPGPU_top.scala 119:24]
  wire [3:0] sm2L2Arb_io_memReqOut_bits_source; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqOut_bits_address; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memReqOut_bits_mask; // @[GPGPU_top.scala 119:24]
  wire [255:0] sm2L2Arb_io_memReqOut_bits_data; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memRspIn_ready; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memRspIn_valid; // @[GPGPU_top.scala 119:24]
  wire [3:0] sm2L2Arb_io_memRspIn_bits_source; // @[GPGPU_top.scala 119:24]
  wire [255:0] sm2L2Arb_io_memRspIn_bits_data; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspIn_bits_address; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memRspVecOut_0_ready; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memRspVecOut_0_valid; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_addr; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_0; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_1; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_2; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_3; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_4; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_5; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_6; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_0_bits_d_data_7; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memRspVecOut_0_bits_d_source; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memRspVecOut_1_ready; // @[GPGPU_top.scala 119:24]
  wire  sm2L2Arb_io_memRspVecOut_1_valid; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_addr; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_0; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_1; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_2; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_3; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_4; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_5; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_6; // @[GPGPU_top.scala 119:24]
  wire [31:0] sm2L2Arb_io_memRspVecOut_1_bits_d_data_7; // @[GPGPU_top.scala 119:24]
  wire [2:0] sm2L2Arb_io_memRspVecOut_1_bits_d_source; // @[GPGPU_top.scala 119:24]
  CTAinterface cta ( // @[GPGPU_top.scala 116:19]
    .clock(cta_clock),
    .reset(cta_reset),
    .io_host2CTA_ready(cta_io_host2CTA_ready),
    .io_host2CTA_valid(cta_io_host2CTA_valid),
    .io_host2CTA_bits_host_wg_id(cta_io_host2CTA_bits_host_wg_id),
    .io_host2CTA_bits_host_num_wf(cta_io_host2CTA_bits_host_num_wf),
    .io_host2CTA_bits_host_wf_size(cta_io_host2CTA_bits_host_wf_size),
    .io_host2CTA_bits_host_start_pc(cta_io_host2CTA_bits_host_start_pc),
    .io_host2CTA_bits_host_vgpr_size_total(cta_io_host2CTA_bits_host_vgpr_size_total),
    .io_host2CTA_bits_host_sgpr_size_total(cta_io_host2CTA_bits_host_sgpr_size_total),
    .io_host2CTA_bits_host_lds_size_total(cta_io_host2CTA_bits_host_lds_size_total),
    .io_host2CTA_bits_host_gds_size_total(cta_io_host2CTA_bits_host_gds_size_total),
    .io_host2CTA_bits_host_vgpr_size_per_wf(cta_io_host2CTA_bits_host_vgpr_size_per_wf),
    .io_host2CTA_bits_host_sgpr_size_per_wf(cta_io_host2CTA_bits_host_sgpr_size_per_wf),
    .io_CTA2host_ready(cta_io_CTA2host_ready),
    .io_CTA2host_valid(cta_io_CTA2host_valid),
    .io_CTA2host_bits_inflight_wg_buffer_host_wf_done_wg_id(cta_io_CTA2host_bits_inflight_wg_buffer_host_wf_done_wg_id),
    .io_CTA2warp_0_ready(cta_io_CTA2warp_0_ready),
    .io_CTA2warp_0_valid(cta_io_CTA2warp_0_valid),
    .io_CTA2warp_0_bits_dispatch2cu_wg_wf_count(cta_io_CTA2warp_0_bits_dispatch2cu_wg_wf_count),
    .io_CTA2warp_0_bits_dispatch2cu_wf_size_dispatch(cta_io_CTA2warp_0_bits_dispatch2cu_wf_size_dispatch),
    .io_CTA2warp_0_bits_dispatch2cu_sgpr_base_dispatch(cta_io_CTA2warp_0_bits_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2warp_0_bits_dispatch2cu_vgpr_base_dispatch(cta_io_CTA2warp_0_bits_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2warp_0_bits_dispatch2cu_wf_tag_dispatch(cta_io_CTA2warp_0_bits_dispatch2cu_wf_tag_dispatch),
    .io_CTA2warp_0_bits_dispatch2cu_lds_base_dispatch(cta_io_CTA2warp_0_bits_dispatch2cu_lds_base_dispatch),
    .io_CTA2warp_0_bits_dispatch2cu_start_pc_dispatch(cta_io_CTA2warp_0_bits_dispatch2cu_start_pc_dispatch),
    .io_CTA2warp_1_ready(cta_io_CTA2warp_1_ready),
    .io_CTA2warp_1_valid(cta_io_CTA2warp_1_valid),
    .io_CTA2warp_1_bits_dispatch2cu_wg_wf_count(cta_io_CTA2warp_1_bits_dispatch2cu_wg_wf_count),
    .io_CTA2warp_1_bits_dispatch2cu_wf_size_dispatch(cta_io_CTA2warp_1_bits_dispatch2cu_wf_size_dispatch),
    .io_CTA2warp_1_bits_dispatch2cu_sgpr_base_dispatch(cta_io_CTA2warp_1_bits_dispatch2cu_sgpr_base_dispatch),
    .io_CTA2warp_1_bits_dispatch2cu_vgpr_base_dispatch(cta_io_CTA2warp_1_bits_dispatch2cu_vgpr_base_dispatch),
    .io_CTA2warp_1_bits_dispatch2cu_wf_tag_dispatch(cta_io_CTA2warp_1_bits_dispatch2cu_wf_tag_dispatch),
    .io_CTA2warp_1_bits_dispatch2cu_lds_base_dispatch(cta_io_CTA2warp_1_bits_dispatch2cu_lds_base_dispatch),
    .io_CTA2warp_1_bits_dispatch2cu_start_pc_dispatch(cta_io_CTA2warp_1_bits_dispatch2cu_start_pc_dispatch),
    .io_warp2CTA_0_valid(cta_io_warp2CTA_0_valid),
    .io_warp2CTA_0_bits_cu2dispatch_wf_tag_done(cta_io_warp2CTA_0_bits_cu2dispatch_wf_tag_done),
    .io_warp2CTA_1_valid(cta_io_warp2CTA_1_valid),
    .io_warp2CTA_1_bits_cu2dispatch_wf_tag_done(cta_io_warp2CTA_1_bits_cu2dispatch_wf_tag_done)
  );
  SM_wrapper SM_wrapper ( // @[GPGPU_top.scala 117:47]
    .clock(SM_wrapper_clock),
    .reset(SM_wrapper_reset),
    .io_CTAreq_ready(SM_wrapper_io_CTAreq_ready),
    .io_CTAreq_valid(SM_wrapper_io_CTAreq_valid),
    .io_CTAreq_bits_dispatch2cu_wg_wf_count(SM_wrapper_io_CTAreq_bits_dispatch2cu_wg_wf_count),
    .io_CTAreq_bits_dispatch2cu_wf_size_dispatch(SM_wrapper_io_CTAreq_bits_dispatch2cu_wf_size_dispatch),
    .io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch(SM_wrapper_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch(SM_wrapper_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_wf_tag_dispatch(SM_wrapper_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch),
    .io_CTAreq_bits_dispatch2cu_lds_base_dispatch(SM_wrapper_io_CTAreq_bits_dispatch2cu_lds_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_start_pc_dispatch(SM_wrapper_io_CTAreq_bits_dispatch2cu_start_pc_dispatch),
    .io_CTArsp_valid(SM_wrapper_io_CTArsp_valid),
    .io_CTArsp_bits_cu2dispatch_wf_tag_done(SM_wrapper_io_CTArsp_bits_cu2dispatch_wf_tag_done),
    .io_memRsp_ready(SM_wrapper_io_memRsp_ready),
    .io_memRsp_valid(SM_wrapper_io_memRsp_valid),
    .io_memRsp_bits_d_addr(SM_wrapper_io_memRsp_bits_d_addr),
    .io_memRsp_bits_d_data_0(SM_wrapper_io_memRsp_bits_d_data_0),
    .io_memRsp_bits_d_data_1(SM_wrapper_io_memRsp_bits_d_data_1),
    .io_memRsp_bits_d_data_2(SM_wrapper_io_memRsp_bits_d_data_2),
    .io_memRsp_bits_d_data_3(SM_wrapper_io_memRsp_bits_d_data_3),
    .io_memRsp_bits_d_data_4(SM_wrapper_io_memRsp_bits_d_data_4),
    .io_memRsp_bits_d_data_5(SM_wrapper_io_memRsp_bits_d_data_5),
    .io_memRsp_bits_d_data_6(SM_wrapper_io_memRsp_bits_d_data_6),
    .io_memRsp_bits_d_data_7(SM_wrapper_io_memRsp_bits_d_data_7),
    .io_memRsp_bits_d_source(SM_wrapper_io_memRsp_bits_d_source),
    .io_memReq_ready(SM_wrapper_io_memReq_ready),
    .io_memReq_valid(SM_wrapper_io_memReq_valid),
    .io_memReq_bits_a_opcode(SM_wrapper_io_memReq_bits_a_opcode),
    .io_memReq_bits_a_addr(SM_wrapper_io_memReq_bits_a_addr),
    .io_memReq_bits_a_data_0(SM_wrapper_io_memReq_bits_a_data_0),
    .io_memReq_bits_a_data_1(SM_wrapper_io_memReq_bits_a_data_1),
    .io_memReq_bits_a_data_2(SM_wrapper_io_memReq_bits_a_data_2),
    .io_memReq_bits_a_data_3(SM_wrapper_io_memReq_bits_a_data_3),
    .io_memReq_bits_a_data_4(SM_wrapper_io_memReq_bits_a_data_4),
    .io_memReq_bits_a_data_5(SM_wrapper_io_memReq_bits_a_data_5),
    .io_memReq_bits_a_data_6(SM_wrapper_io_memReq_bits_a_data_6),
    .io_memReq_bits_a_data_7(SM_wrapper_io_memReq_bits_a_data_7),
    .io_memReq_bits_a_mask_0(SM_wrapper_io_memReq_bits_a_mask_0),
    .io_memReq_bits_a_mask_1(SM_wrapper_io_memReq_bits_a_mask_1),
    .io_memReq_bits_a_mask_2(SM_wrapper_io_memReq_bits_a_mask_2),
    .io_memReq_bits_a_mask_3(SM_wrapper_io_memReq_bits_a_mask_3),
    .io_memReq_bits_a_mask_4(SM_wrapper_io_memReq_bits_a_mask_4),
    .io_memReq_bits_a_mask_5(SM_wrapper_io_memReq_bits_a_mask_5),
    .io_memReq_bits_a_mask_6(SM_wrapper_io_memReq_bits_a_mask_6),
    .io_memReq_bits_a_mask_7(SM_wrapper_io_memReq_bits_a_mask_7),
    .io_memReq_bits_a_source(SM_wrapper_io_memReq_bits_a_source)
  );
  SM_wrapper SM_wrapper_1 ( // @[GPGPU_top.scala 117:47]
    .clock(SM_wrapper_1_clock),
    .reset(SM_wrapper_1_reset),
    .io_CTAreq_ready(SM_wrapper_1_io_CTAreq_ready),
    .io_CTAreq_valid(SM_wrapper_1_io_CTAreq_valid),
    .io_CTAreq_bits_dispatch2cu_wg_wf_count(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wg_wf_count),
    .io_CTAreq_bits_dispatch2cu_wf_size_dispatch(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wf_size_dispatch),
    .io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_wf_tag_dispatch(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch),
    .io_CTAreq_bits_dispatch2cu_lds_base_dispatch(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_lds_base_dispatch),
    .io_CTAreq_bits_dispatch2cu_start_pc_dispatch(SM_wrapper_1_io_CTAreq_bits_dispatch2cu_start_pc_dispatch),
    .io_CTArsp_valid(SM_wrapper_1_io_CTArsp_valid),
    .io_CTArsp_bits_cu2dispatch_wf_tag_done(SM_wrapper_1_io_CTArsp_bits_cu2dispatch_wf_tag_done),
    .io_memRsp_ready(SM_wrapper_1_io_memRsp_ready),
    .io_memRsp_valid(SM_wrapper_1_io_memRsp_valid),
    .io_memRsp_bits_d_addr(SM_wrapper_1_io_memRsp_bits_d_addr),
    .io_memRsp_bits_d_data_0(SM_wrapper_1_io_memRsp_bits_d_data_0),
    .io_memRsp_bits_d_data_1(SM_wrapper_1_io_memRsp_bits_d_data_1),
    .io_memRsp_bits_d_data_2(SM_wrapper_1_io_memRsp_bits_d_data_2),
    .io_memRsp_bits_d_data_3(SM_wrapper_1_io_memRsp_bits_d_data_3),
    .io_memRsp_bits_d_data_4(SM_wrapper_1_io_memRsp_bits_d_data_4),
    .io_memRsp_bits_d_data_5(SM_wrapper_1_io_memRsp_bits_d_data_5),
    .io_memRsp_bits_d_data_6(SM_wrapper_1_io_memRsp_bits_d_data_6),
    .io_memRsp_bits_d_data_7(SM_wrapper_1_io_memRsp_bits_d_data_7),
    .io_memRsp_bits_d_source(SM_wrapper_1_io_memRsp_bits_d_source),
    .io_memReq_ready(SM_wrapper_1_io_memReq_ready),
    .io_memReq_valid(SM_wrapper_1_io_memReq_valid),
    .io_memReq_bits_a_opcode(SM_wrapper_1_io_memReq_bits_a_opcode),
    .io_memReq_bits_a_addr(SM_wrapper_1_io_memReq_bits_a_addr),
    .io_memReq_bits_a_data_0(SM_wrapper_1_io_memReq_bits_a_data_0),
    .io_memReq_bits_a_data_1(SM_wrapper_1_io_memReq_bits_a_data_1),
    .io_memReq_bits_a_data_2(SM_wrapper_1_io_memReq_bits_a_data_2),
    .io_memReq_bits_a_data_3(SM_wrapper_1_io_memReq_bits_a_data_3),
    .io_memReq_bits_a_data_4(SM_wrapper_1_io_memReq_bits_a_data_4),
    .io_memReq_bits_a_data_5(SM_wrapper_1_io_memReq_bits_a_data_5),
    .io_memReq_bits_a_data_6(SM_wrapper_1_io_memReq_bits_a_data_6),
    .io_memReq_bits_a_data_7(SM_wrapper_1_io_memReq_bits_a_data_7),
    .io_memReq_bits_a_mask_0(SM_wrapper_1_io_memReq_bits_a_mask_0),
    .io_memReq_bits_a_mask_1(SM_wrapper_1_io_memReq_bits_a_mask_1),
    .io_memReq_bits_a_mask_2(SM_wrapper_1_io_memReq_bits_a_mask_2),
    .io_memReq_bits_a_mask_3(SM_wrapper_1_io_memReq_bits_a_mask_3),
    .io_memReq_bits_a_mask_4(SM_wrapper_1_io_memReq_bits_a_mask_4),
    .io_memReq_bits_a_mask_5(SM_wrapper_1_io_memReq_bits_a_mask_5),
    .io_memReq_bits_a_mask_6(SM_wrapper_1_io_memReq_bits_a_mask_6),
    .io_memReq_bits_a_mask_7(SM_wrapper_1_io_memReq_bits_a_mask_7),
    .io_memReq_bits_a_source(SM_wrapper_1_io_memReq_bits_a_source)
  );
  Scheduler l2cache ( // @[GPGPU_top.scala 118:21]
    .clock(l2cache_clock),
    .reset(l2cache_reset),
    .io_in_a_ready(l2cache_io_in_a_ready),
    .io_in_a_valid(l2cache_io_in_a_valid),
    .io_in_a_bits_opcode(l2cache_io_in_a_bits_opcode),
    .io_in_a_bits_source(l2cache_io_in_a_bits_source),
    .io_in_a_bits_address(l2cache_io_in_a_bits_address),
    .io_in_a_bits_mask(l2cache_io_in_a_bits_mask),
    .io_in_a_bits_data(l2cache_io_in_a_bits_data),
    .io_in_d_ready(l2cache_io_in_d_ready),
    .io_in_d_valid(l2cache_io_in_d_valid),
    .io_in_d_bits_source(l2cache_io_in_d_bits_source),
    .io_in_d_bits_data(l2cache_io_in_d_bits_data),
    .io_in_d_bits_address(l2cache_io_in_d_bits_address),
    .io_out_a_ready(l2cache_io_out_a_ready),
    .io_out_a_valid(l2cache_io_out_a_valid),
    .io_out_a_bits_opcode(l2cache_io_out_a_bits_opcode),
    .io_out_a_bits_source(l2cache_io_out_a_bits_source),
    .io_out_a_bits_address(l2cache_io_out_a_bits_address),
    .io_out_a_bits_mask(l2cache_io_out_a_bits_mask),
    .io_out_a_bits_data(l2cache_io_out_a_bits_data),
    .io_out_d_ready(l2cache_io_out_d_ready),
    .io_out_d_valid(l2cache_io_out_d_valid),
    .io_out_d_bits_opcode(l2cache_io_out_d_bits_opcode),
    .io_out_d_bits_source(l2cache_io_out_d_bits_source),
    .io_out_d_bits_data(l2cache_io_out_d_bits_data)
  );
  SM2L2Arbiter sm2L2Arb ( // @[GPGPU_top.scala 119:24]
    .io_memReqVecIn_0_ready(sm2L2Arb_io_memReqVecIn_0_ready),
    .io_memReqVecIn_0_valid(sm2L2Arb_io_memReqVecIn_0_valid),
    .io_memReqVecIn_0_bits_a_opcode(sm2L2Arb_io_memReqVecIn_0_bits_a_opcode),
    .io_memReqVecIn_0_bits_a_addr(sm2L2Arb_io_memReqVecIn_0_bits_a_addr),
    .io_memReqVecIn_0_bits_a_data_0(sm2L2Arb_io_memReqVecIn_0_bits_a_data_0),
    .io_memReqVecIn_0_bits_a_data_1(sm2L2Arb_io_memReqVecIn_0_bits_a_data_1),
    .io_memReqVecIn_0_bits_a_data_2(sm2L2Arb_io_memReqVecIn_0_bits_a_data_2),
    .io_memReqVecIn_0_bits_a_data_3(sm2L2Arb_io_memReqVecIn_0_bits_a_data_3),
    .io_memReqVecIn_0_bits_a_data_4(sm2L2Arb_io_memReqVecIn_0_bits_a_data_4),
    .io_memReqVecIn_0_bits_a_data_5(sm2L2Arb_io_memReqVecIn_0_bits_a_data_5),
    .io_memReqVecIn_0_bits_a_data_6(sm2L2Arb_io_memReqVecIn_0_bits_a_data_6),
    .io_memReqVecIn_0_bits_a_data_7(sm2L2Arb_io_memReqVecIn_0_bits_a_data_7),
    .io_memReqVecIn_0_bits_a_mask_0(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_0),
    .io_memReqVecIn_0_bits_a_mask_1(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_1),
    .io_memReqVecIn_0_bits_a_mask_2(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_2),
    .io_memReqVecIn_0_bits_a_mask_3(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_3),
    .io_memReqVecIn_0_bits_a_mask_4(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_4),
    .io_memReqVecIn_0_bits_a_mask_5(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_5),
    .io_memReqVecIn_0_bits_a_mask_6(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_6),
    .io_memReqVecIn_0_bits_a_mask_7(sm2L2Arb_io_memReqVecIn_0_bits_a_mask_7),
    .io_memReqVecIn_0_bits_a_source(sm2L2Arb_io_memReqVecIn_0_bits_a_source),
    .io_memReqVecIn_1_ready(sm2L2Arb_io_memReqVecIn_1_ready),
    .io_memReqVecIn_1_valid(sm2L2Arb_io_memReqVecIn_1_valid),
    .io_memReqVecIn_1_bits_a_opcode(sm2L2Arb_io_memReqVecIn_1_bits_a_opcode),
    .io_memReqVecIn_1_bits_a_addr(sm2L2Arb_io_memReqVecIn_1_bits_a_addr),
    .io_memReqVecIn_1_bits_a_data_0(sm2L2Arb_io_memReqVecIn_1_bits_a_data_0),
    .io_memReqVecIn_1_bits_a_data_1(sm2L2Arb_io_memReqVecIn_1_bits_a_data_1),
    .io_memReqVecIn_1_bits_a_data_2(sm2L2Arb_io_memReqVecIn_1_bits_a_data_2),
    .io_memReqVecIn_1_bits_a_data_3(sm2L2Arb_io_memReqVecIn_1_bits_a_data_3),
    .io_memReqVecIn_1_bits_a_data_4(sm2L2Arb_io_memReqVecIn_1_bits_a_data_4),
    .io_memReqVecIn_1_bits_a_data_5(sm2L2Arb_io_memReqVecIn_1_bits_a_data_5),
    .io_memReqVecIn_1_bits_a_data_6(sm2L2Arb_io_memReqVecIn_1_bits_a_data_6),
    .io_memReqVecIn_1_bits_a_data_7(sm2L2Arb_io_memReqVecIn_1_bits_a_data_7),
    .io_memReqVecIn_1_bits_a_mask_0(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_0),
    .io_memReqVecIn_1_bits_a_mask_1(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_1),
    .io_memReqVecIn_1_bits_a_mask_2(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_2),
    .io_memReqVecIn_1_bits_a_mask_3(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_3),
    .io_memReqVecIn_1_bits_a_mask_4(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_4),
    .io_memReqVecIn_1_bits_a_mask_5(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_5),
    .io_memReqVecIn_1_bits_a_mask_6(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_6),
    .io_memReqVecIn_1_bits_a_mask_7(sm2L2Arb_io_memReqVecIn_1_bits_a_mask_7),
    .io_memReqVecIn_1_bits_a_source(sm2L2Arb_io_memReqVecIn_1_bits_a_source),
    .io_memReqOut_ready(sm2L2Arb_io_memReqOut_ready),
    .io_memReqOut_valid(sm2L2Arb_io_memReqOut_valid),
    .io_memReqOut_bits_opcode(sm2L2Arb_io_memReqOut_bits_opcode),
    .io_memReqOut_bits_source(sm2L2Arb_io_memReqOut_bits_source),
    .io_memReqOut_bits_address(sm2L2Arb_io_memReqOut_bits_address),
    .io_memReqOut_bits_mask(sm2L2Arb_io_memReqOut_bits_mask),
    .io_memReqOut_bits_data(sm2L2Arb_io_memReqOut_bits_data),
    .io_memRspIn_ready(sm2L2Arb_io_memRspIn_ready),
    .io_memRspIn_valid(sm2L2Arb_io_memRspIn_valid),
    .io_memRspIn_bits_source(sm2L2Arb_io_memRspIn_bits_source),
    .io_memRspIn_bits_data(sm2L2Arb_io_memRspIn_bits_data),
    .io_memRspIn_bits_address(sm2L2Arb_io_memRspIn_bits_address),
    .io_memRspVecOut_0_ready(sm2L2Arb_io_memRspVecOut_0_ready),
    .io_memRspVecOut_0_valid(sm2L2Arb_io_memRspVecOut_0_valid),
    .io_memRspVecOut_0_bits_d_addr(sm2L2Arb_io_memRspVecOut_0_bits_d_addr),
    .io_memRspVecOut_0_bits_d_data_0(sm2L2Arb_io_memRspVecOut_0_bits_d_data_0),
    .io_memRspVecOut_0_bits_d_data_1(sm2L2Arb_io_memRspVecOut_0_bits_d_data_1),
    .io_memRspVecOut_0_bits_d_data_2(sm2L2Arb_io_memRspVecOut_0_bits_d_data_2),
    .io_memRspVecOut_0_bits_d_data_3(sm2L2Arb_io_memRspVecOut_0_bits_d_data_3),
    .io_memRspVecOut_0_bits_d_data_4(sm2L2Arb_io_memRspVecOut_0_bits_d_data_4),
    .io_memRspVecOut_0_bits_d_data_5(sm2L2Arb_io_memRspVecOut_0_bits_d_data_5),
    .io_memRspVecOut_0_bits_d_data_6(sm2L2Arb_io_memRspVecOut_0_bits_d_data_6),
    .io_memRspVecOut_0_bits_d_data_7(sm2L2Arb_io_memRspVecOut_0_bits_d_data_7),
    .io_memRspVecOut_0_bits_d_source(sm2L2Arb_io_memRspVecOut_0_bits_d_source),
    .io_memRspVecOut_1_ready(sm2L2Arb_io_memRspVecOut_1_ready),
    .io_memRspVecOut_1_valid(sm2L2Arb_io_memRspVecOut_1_valid),
    .io_memRspVecOut_1_bits_d_addr(sm2L2Arb_io_memRspVecOut_1_bits_d_addr),
    .io_memRspVecOut_1_bits_d_data_0(sm2L2Arb_io_memRspVecOut_1_bits_d_data_0),
    .io_memRspVecOut_1_bits_d_data_1(sm2L2Arb_io_memRspVecOut_1_bits_d_data_1),
    .io_memRspVecOut_1_bits_d_data_2(sm2L2Arb_io_memRspVecOut_1_bits_d_data_2),
    .io_memRspVecOut_1_bits_d_data_3(sm2L2Arb_io_memRspVecOut_1_bits_d_data_3),
    .io_memRspVecOut_1_bits_d_data_4(sm2L2Arb_io_memRspVecOut_1_bits_d_data_4),
    .io_memRspVecOut_1_bits_d_data_5(sm2L2Arb_io_memRspVecOut_1_bits_d_data_5),
    .io_memRspVecOut_1_bits_d_data_6(sm2L2Arb_io_memRspVecOut_1_bits_d_data_6),
    .io_memRspVecOut_1_bits_d_data_7(sm2L2Arb_io_memRspVecOut_1_bits_d_data_7),
    .io_memRspVecOut_1_bits_d_source(sm2L2Arb_io_memRspVecOut_1_bits_d_source)
  );
  assign io_host_req_ready = cta_io_host2CTA_ready; // @[GPGPU_top.scala 133:14]
  assign io_host_rsp_valid = cta_io_CTA2host_valid; // @[GPGPU_top.scala 132:14]
  assign io_host_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id =
    cta_io_CTA2host_bits_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 132:14]
  assign io_out_a_valid = l2cache_io_out_a_valid; // @[GPGPU_top.scala 129:20]
  assign io_out_a_bits_opcode = l2cache_io_out_a_bits_opcode; // @[GPGPU_top.scala 129:20]
  assign io_out_a_bits_source = l2cache_io_out_a_bits_source; // @[GPGPU_top.scala 129:20]
  assign io_out_a_bits_address = l2cache_io_out_a_bits_address; // @[GPGPU_top.scala 129:20]
  assign io_out_a_bits_mask = l2cache_io_out_a_bits_mask; // @[GPGPU_top.scala 129:20]
  assign io_out_a_bits_data = l2cache_io_out_a_bits_data; // @[GPGPU_top.scala 129:20]
  assign io_out_d_ready = l2cache_io_out_d_ready; // @[GPGPU_top.scala 130:20]
  assign cta_clock = clock;
  assign cta_reset = reset;
  assign cta_io_host2CTA_valid = io_host_req_valid; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_wg_id = io_host_req_bits_host_wg_id; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_num_wf = io_host_req_bits_host_num_wf; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_wf_size = io_host_req_bits_host_wf_size; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_start_pc = io_host_req_bits_host_start_pc; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_vgpr_size_total = io_host_req_bits_host_vgpr_size_total; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_sgpr_size_total = io_host_req_bits_host_sgpr_size_total; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_lds_size_total = io_host_req_bits_host_lds_size_total; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_gds_size_total = io_host_req_bits_host_gds_size_total; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_vgpr_size_per_wf = io_host_req_bits_host_vgpr_size_per_wf; // @[GPGPU_top.scala 133:14]
  assign cta_io_host2CTA_bits_host_sgpr_size_per_wf = io_host_req_bits_host_sgpr_size_per_wf; // @[GPGPU_top.scala 133:14]
  assign cta_io_CTA2host_ready = io_host_rsp_ready; // @[GPGPU_top.scala 132:14]
  assign cta_io_CTA2warp_0_ready = SM_wrapper_io_CTAreq_ready; // @[GPGPU_top.scala 117:{25,25}]
  assign cta_io_CTA2warp_1_ready = SM_wrapper_1_io_CTAreq_ready; // @[GPGPU_top.scala 117:{25,25}]
  assign cta_io_warp2CTA_0_valid = SM_wrapper_io_CTArsp_valid; // @[GPGPU_top.scala 117:{25,25}]
  assign cta_io_warp2CTA_0_bits_cu2dispatch_wf_tag_done = SM_wrapper_io_CTArsp_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 117:{25,25}]
  assign cta_io_warp2CTA_1_valid = SM_wrapper_1_io_CTArsp_valid; // @[GPGPU_top.scala 117:{25,25}]
  assign cta_io_warp2CTA_1_bits_cu2dispatch_wf_tag_done = SM_wrapper_1_io_CTArsp_bits_cu2dispatch_wf_tag_done; // @[GPGPU_top.scala 117:{25,25}]
  assign SM_wrapper_clock = clock;
  assign SM_wrapper_reset = reset;
  assign SM_wrapper_io_CTAreq_valid = cta_io_CTA2warp_0_valid; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_wg_wf_count = cta_io_CTA2warp_0_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_wf_size_dispatch = cta_io_CTA2warp_0_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch =
    cta_io_CTA2warp_0_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch =
    cta_io_CTA2warp_0_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch = cta_io_CTA2warp_0_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_lds_base_dispatch = cta_io_CTA2warp_0_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_CTAreq_bits_dispatch2cu_start_pc_dispatch = cta_io_CTA2warp_0_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_io_memRsp_valid = sm2L2Arb_io_memRspVecOut_0_valid; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_addr = sm2L2Arb_io_memRspVecOut_0_bits_d_addr; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_0 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_0; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_1 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_1; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_2 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_2; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_3 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_3; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_4 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_4; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_5 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_5; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_6 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_6; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_data_7 = sm2L2Arb_io_memRspVecOut_0_bits_d_data_7; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memRsp_bits_d_source = sm2L2Arb_io_memRspVecOut_0_bits_d_source; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_io_memReq_ready = sm2L2Arb_io_memReqVecIn_0_ready; // @[GPGPU_top.scala 117:25 125:32]
  assign SM_wrapper_1_clock = clock;
  assign SM_wrapper_1_reset = reset;
  assign SM_wrapper_1_io_CTAreq_valid = cta_io_CTA2warp_1_valid; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wg_wf_count = cta_io_CTA2warp_1_bits_dispatch2cu_wg_wf_count; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wf_size_dispatch = cta_io_CTA2warp_1_bits_dispatch2cu_wf_size_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_sgpr_base_dispatch =
    cta_io_CTA2warp_1_bits_dispatch2cu_sgpr_base_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_vgpr_base_dispatch =
    cta_io_CTA2warp_1_bits_dispatch2cu_vgpr_base_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_wf_tag_dispatch = cta_io_CTA2warp_1_bits_dispatch2cu_wf_tag_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_lds_base_dispatch =
    cta_io_CTA2warp_1_bits_dispatch2cu_lds_base_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_CTAreq_bits_dispatch2cu_start_pc_dispatch =
    cta_io_CTA2warp_1_bits_dispatch2cu_start_pc_dispatch; // @[GPGPU_top.scala 117:25 122:23]
  assign SM_wrapper_1_io_memRsp_valid = sm2L2Arb_io_memRspVecOut_1_valid; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_addr = sm2L2Arb_io_memRspVecOut_1_bits_d_addr; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_0 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_0; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_1 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_1; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_2 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_2; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_3 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_3; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_4 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_4; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_5 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_5; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_6 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_6; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_data_7 = sm2L2Arb_io_memRspVecOut_1_bits_d_data_7; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memRsp_bits_d_source = sm2L2Arb_io_memRspVecOut_1_bits_d_source; // @[GPGPU_top.scala 117:25 124:26]
  assign SM_wrapper_1_io_memReq_ready = sm2L2Arb_io_memReqVecIn_1_ready; // @[GPGPU_top.scala 117:25 125:32]
  assign l2cache_clock = clock;
  assign l2cache_reset = reset;
  assign l2cache_io_in_a_valid = sm2L2Arb_io_memReqOut_valid; // @[GPGPU_top.scala 128:19]
  assign l2cache_io_in_a_bits_opcode = sm2L2Arb_io_memReqOut_bits_opcode; // @[GPGPU_top.scala 128:19]
  assign l2cache_io_in_a_bits_source = sm2L2Arb_io_memReqOut_bits_source; // @[GPGPU_top.scala 128:19]
  assign l2cache_io_in_a_bits_address = sm2L2Arb_io_memReqOut_bits_address; // @[GPGPU_top.scala 128:19]
  assign l2cache_io_in_a_bits_mask = sm2L2Arb_io_memReqOut_bits_mask; // @[GPGPU_top.scala 128:19]
  assign l2cache_io_in_a_bits_data = sm2L2Arb_io_memReqOut_bits_data; // @[GPGPU_top.scala 128:19]
  assign l2cache_io_in_d_ready = sm2L2Arb_io_memRspIn_ready; // @[GPGPU_top.scala 131:24]
  assign l2cache_io_out_a_ready = io_out_a_ready; // @[GPGPU_top.scala 129:20]
  assign l2cache_io_out_d_valid = io_out_d_valid; // @[GPGPU_top.scala 130:20]
  assign l2cache_io_out_d_bits_opcode = io_out_d_bits_opcode; // @[GPGPU_top.scala 130:20]
  assign l2cache_io_out_d_bits_source = io_out_d_bits_source; // @[GPGPU_top.scala 130:20]
  assign l2cache_io_out_d_bits_data = io_out_d_bits_data; // @[GPGPU_top.scala 130:20]
  assign sm2L2Arb_io_memReqVecIn_0_valid = SM_wrapper_io_memReq_valid; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_opcode = SM_wrapper_io_memReq_bits_a_opcode; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_addr = SM_wrapper_io_memReq_bits_a_addr; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_0 = SM_wrapper_io_memReq_bits_a_data_0; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_1 = SM_wrapper_io_memReq_bits_a_data_1; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_2 = SM_wrapper_io_memReq_bits_a_data_2; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_3 = SM_wrapper_io_memReq_bits_a_data_3; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_4 = SM_wrapper_io_memReq_bits_a_data_4; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_5 = SM_wrapper_io_memReq_bits_a_data_5; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_6 = SM_wrapper_io_memReq_bits_a_data_6; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_data_7 = SM_wrapper_io_memReq_bits_a_data_7; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_0 = SM_wrapper_io_memReq_bits_a_mask_0; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_1 = SM_wrapper_io_memReq_bits_a_mask_1; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_2 = SM_wrapper_io_memReq_bits_a_mask_2; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_3 = SM_wrapper_io_memReq_bits_a_mask_3; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_4 = SM_wrapper_io_memReq_bits_a_mask_4; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_5 = SM_wrapper_io_memReq_bits_a_mask_5; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_6 = SM_wrapper_io_memReq_bits_a_mask_6; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_mask_7 = SM_wrapper_io_memReq_bits_a_mask_7; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_0_bits_a_source = SM_wrapper_io_memReq_bits_a_source; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_valid = SM_wrapper_1_io_memReq_valid; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_opcode = SM_wrapper_1_io_memReq_bits_a_opcode; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_addr = SM_wrapper_1_io_memReq_bits_a_addr; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_0 = SM_wrapper_1_io_memReq_bits_a_data_0; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_1 = SM_wrapper_1_io_memReq_bits_a_data_1; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_2 = SM_wrapper_1_io_memReq_bits_a_data_2; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_3 = SM_wrapper_1_io_memReq_bits_a_data_3; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_4 = SM_wrapper_1_io_memReq_bits_a_data_4; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_5 = SM_wrapper_1_io_memReq_bits_a_data_5; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_6 = SM_wrapper_1_io_memReq_bits_a_data_6; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_data_7 = SM_wrapper_1_io_memReq_bits_a_data_7; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_0 = SM_wrapper_1_io_memReq_bits_a_mask_0; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_1 = SM_wrapper_1_io_memReq_bits_a_mask_1; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_2 = SM_wrapper_1_io_memReq_bits_a_mask_2; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_3 = SM_wrapper_1_io_memReq_bits_a_mask_3; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_4 = SM_wrapper_1_io_memReq_bits_a_mask_4; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_5 = SM_wrapper_1_io_memReq_bits_a_mask_5; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_6 = SM_wrapper_1_io_memReq_bits_a_mask_6; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_mask_7 = SM_wrapper_1_io_memReq_bits_a_mask_7; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqVecIn_1_bits_a_source = SM_wrapper_1_io_memReq_bits_a_source; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memReqOut_ready = l2cache_io_in_a_ready; // @[GPGPU_top.scala 128:19]
  assign sm2L2Arb_io_memRspIn_valid = l2cache_io_in_d_valid; // @[GPGPU_top.scala 131:24]
  assign sm2L2Arb_io_memRspIn_bits_source = l2cache_io_in_d_bits_source; // @[GPGPU_top.scala 131:24]
  assign sm2L2Arb_io_memRspIn_bits_data = l2cache_io_in_d_bits_data; // @[GPGPU_top.scala 131:24]
  assign sm2L2Arb_io_memRspIn_bits_address = l2cache_io_in_d_bits_address; // @[GPGPU_top.scala 131:24]
  assign sm2L2Arb_io_memRspVecOut_0_ready = SM_wrapper_io_memRsp_ready; // @[GPGPU_top.scala 117:{25,25}]
  assign sm2L2Arb_io_memRspVecOut_1_ready = SM_wrapper_1_io_memRsp_ready; // @[GPGPU_top.scala 117:{25,25}]
endmodule
module AXI4Lite2CTA(
  input         clock,
  input         reset,
  input  [31:0] io_ctl_aw_awaddr,
  input         io_ctl_aw_awvalid,
  output        io_ctl_aw_awready,
  input  [11:0] io_ctl_aw_awid,
  input  [31:0] io_ctl_w_wdata,
  input         io_ctl_w_wvalid,
  output        io_ctl_w_wready,
  output        io_ctl_b_bvalid,
  input         io_ctl_b_bready,
  output [11:0] io_ctl_b_bid,
  input  [31:0] io_ctl_ar_araddr,
  input         io_ctl_ar_arvalid,
  output        io_ctl_ar_arready,
  input  [11:0] io_ctl_ar_arid,
  output [31:0] io_ctl_r_rdata,
  output        io_ctl_r_rvalid,
  input         io_ctl_r_rready,
  output [11:0] io_ctl_r_rid,
  input         io_data_ready,
  output        io_data_valid,
  output [4:0]  io_data_bits_host_wg_id,
  output [2:0]  io_data_bits_host_num_wf,
  output [9:0]  io_data_bits_host_wf_size,
  output [31:0] io_data_bits_host_start_pc,
  output [12:0] io_data_bits_host_vgpr_size_total,
  output [12:0] io_data_bits_host_sgpr_size_total,
  output [12:0] io_data_bits_host_lds_size_total,
  output [10:0] io_data_bits_host_gds_size_total,
  output [12:0] io_data_bits_host_vgpr_size_per_wf,
  output [12:0] io_data_bits_host_sgpr_size_per_wf,
  output        io_rsp_ready,
  input         io_rsp_valid,
  input  [4:0]  io_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_1; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_2; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_3; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_4; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_5; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_6; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_7; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_8; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_9; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_10; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_11; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_12; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_13; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_14; // @[AXI4Lite2CTA.scala 50:21]
  reg [31:0] regs_15; // @[AXI4Lite2CTA.scala 50:21]
  wire [31:0] _GEN_1 = io_rsp_valid & ~regs_15[0] ? 32'h1 : regs_15; // @[AXI4Lite2CTA.scala 53:35 55:13 50:21]
  wire [31:0] _GEN_2 = io_rsp_valid & ~regs_15[0] ? {{27'd0}, io_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id} :
    regs_14; // @[AXI4Lite2CTA.scala 53:35 56:13 50:21]
  reg [2:0] state; // @[AXI4Lite2CTA.scala 60:22]
  reg  awready; // @[AXI4Lite2CTA.scala 62:24]
  reg  wready; // @[AXI4Lite2CTA.scala 63:23]
  reg  bvalid; // @[AXI4Lite2CTA.scala 64:23]
  reg  arready; // @[AXI4Lite2CTA.scala 67:24]
  reg  rvalid; // @[AXI4Lite2CTA.scala 68:23]
  reg [31:0] addr; // @[AXI4Lite2CTA.scala 71:21]
  reg  write; // @[AXI4Lite2CTA.scala 74:22]
  reg [31:0] dataOut; // @[AXI4Lite2CTA.scala 75:24]
  reg [11:0] transaction_id; // @[AXI4Lite2CTA.scala 77:31]
  wire [31:0] _GEN_4 = 4'h1 == addr[3:0] ? regs_1 : regs_0; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_5 = 4'h2 == addr[3:0] ? regs_2 : _GEN_4; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_6 = 4'h3 == addr[3:0] ? regs_3 : _GEN_5; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_7 = 4'h4 == addr[3:0] ? regs_4 : _GEN_6; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_8 = 4'h5 == addr[3:0] ? regs_5 : _GEN_7; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_9 = 4'h6 == addr[3:0] ? regs_6 : _GEN_8; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_10 = 4'h7 == addr[3:0] ? regs_7 : _GEN_9; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_11 = 4'h8 == addr[3:0] ? regs_8 : _GEN_10; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_12 = 4'h9 == addr[3:0] ? regs_9 : _GEN_11; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_13 = 4'ha == addr[3:0] ? regs_10 : _GEN_12; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_14 = 4'hb == addr[3:0] ? regs_11 : _GEN_13; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_15 = 4'hc == addr[3:0] ? regs_12 : _GEN_14; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_16 = 4'hd == addr[3:0] ? regs_13 : _GEN_15; // @[AXI4Lite2CTA.scala 79:{18,18}]
  wire [31:0] _GEN_17 = 4'he == addr[3:0] ? regs_14 : _GEN_16; // @[AXI4Lite2CTA.scala 79:{18,18}]
  reg  out_state; // @[AXI4Lite2CTA.scala 95:24]
  wire  input_valid = regs_0[0]; // @[AXI4Lite2CTA.scala 96:26]
  wire  _T_3 = ~out_state; // @[AXI4Lite2CTA.scala 110:21]
  wire  _GEN_19 = input_valid | out_state; // @[AXI4Lite2CTA.scala 112:25 113:19 95:24]
  wire  _T_5 = io_data_ready & io_data_valid; // @[Decoupled.scala 50:35]
  wire [31:0] _GEN_21 = _T_5 ? 32'h0 : regs_0; // @[AXI4Lite2CTA.scala 117:26 119:16 50:21]
  wire [31:0] _GEN_23 = out_state ? _GEN_21 : regs_0; // @[AXI4Lite2CTA.scala 110:21 50:21]
  wire [31:0] _GEN_25 = ~out_state ? regs_0 : _GEN_23; // @[AXI4Lite2CTA.scala 110:21 50:21]
  wire [2:0] _GEN_66 = io_ctl_r_rready & rvalid ? 3'h0 : state; // @[AXI4Lite2CTA.scala 154:38 155:15 60:22]
  wire  _GEN_67 = io_ctl_r_rready & rvalid ? 1'h0 : 1'h1; // @[AXI4Lite2CTA.scala 153:14 154:38 156:16]
  wire [31:0] _GEN_68 = io_ctl_aw_awvalid & awready ? {{2'd0}, io_ctl_aw_awaddr[31:2]} : addr; // @[AXI4Lite2CTA.scala 161:41 162:14 71:21]
  wire [2:0] _GEN_69 = io_ctl_aw_awvalid & awready ? 3'h4 : state; // @[AXI4Lite2CTA.scala 161:41 163:15 60:22]
  wire  _GEN_70 = io_ctl_aw_awvalid & awready ? 1'h0 : 1'h1; // @[AXI4Lite2CTA.scala 160:15 161:41 164:17]
  wire [2:0] _GEN_71 = io_ctl_w_wvalid & wready ? 3'h5 : state; // @[AXI4Lite2CTA.scala 169:38 170:15 60:22]
  wire [31:0] _GEN_72 = io_ctl_w_wvalid & wready ? io_ctl_w_wdata : dataOut; // @[AXI4Lite2CTA.scala 169:38 171:17 75:24]
  wire  _GEN_73 = io_ctl_w_wvalid & wready | write; // @[AXI4Lite2CTA.scala 169:38 172:15 74:22]
  wire  _GEN_74 = io_ctl_w_wvalid & wready ? 1'h0 : 1'h1; // @[AXI4Lite2CTA.scala 168:14 169:38 173:16]
  wire [2:0] _GEN_75 = io_ctl_b_bready & bvalid ? 3'h0 : state; // @[AXI4Lite2CTA.scala 179:38 180:15 60:22]
  wire  _GEN_76 = io_ctl_b_bready & bvalid ? 1'h0 : 1'h1; // @[AXI4Lite2CTA.scala 178:14 179:38 181:16]
  wire  _GEN_77 = 3'h5 == state ? 1'h0 : wready; // @[AXI4Lite2CTA.scala 127:16 177:14 63:23]
  wire  _GEN_78 = 3'h5 == state ? _GEN_76 : bvalid; // @[AXI4Lite2CTA.scala 127:16 64:23]
  wire [2:0] _GEN_79 = 3'h5 == state ? _GEN_75 : state; // @[AXI4Lite2CTA.scala 127:16 60:22]
  wire  _GEN_80 = 3'h4 == state ? _GEN_74 : _GEN_77; // @[AXI4Lite2CTA.scala 127:16]
  wire [2:0] _GEN_81 = 3'h4 == state ? _GEN_71 : _GEN_79; // @[AXI4Lite2CTA.scala 127:16]
  wire [31:0] _GEN_82 = 3'h4 == state ? _GEN_72 : dataOut; // @[AXI4Lite2CTA.scala 127:16 75:24]
  wire  _GEN_83 = 3'h4 == state ? _GEN_73 : write; // @[AXI4Lite2CTA.scala 127:16 74:22]
  wire  _GEN_84 = 3'h4 == state ? bvalid : _GEN_78; // @[AXI4Lite2CTA.scala 127:16 64:23]
  wire  _GEN_85 = 3'h3 == state ? _GEN_70 : awready; // @[AXI4Lite2CTA.scala 127:16 62:24]
  wire [31:0] _GEN_86 = 3'h3 == state ? _GEN_68 : addr; // @[AXI4Lite2CTA.scala 127:16 71:21]
  wire [2:0] _GEN_87 = 3'h3 == state ? _GEN_69 : _GEN_81; // @[AXI4Lite2CTA.scala 127:16]
  wire  _GEN_88 = 3'h3 == state ? wready : _GEN_80; // @[AXI4Lite2CTA.scala 127:16 63:23]
  wire [31:0] _GEN_89 = 3'h3 == state ? dataOut : _GEN_82; // @[AXI4Lite2CTA.scala 127:16 75:24]
  wire  _GEN_90 = 3'h3 == state ? write : _GEN_83; // @[AXI4Lite2CTA.scala 127:16 74:22]
  wire  _GEN_91 = 3'h3 == state ? bvalid : _GEN_84; // @[AXI4Lite2CTA.scala 127:16 64:23]
  assign io_ctl_aw_awready = awready; // @[AXI4Lite2CTA.scala 83:21]
  assign io_ctl_w_wready = wready; // @[AXI4Lite2CTA.scala 84:19]
  assign io_ctl_b_bvalid = bvalid; // @[AXI4Lite2CTA.scala 85:19]
  assign io_ctl_b_bid = transaction_id; // @[AXI4Lite2CTA.scala 87:16]
  assign io_ctl_ar_arready = arready; // @[AXI4Lite2CTA.scala 89:21]
  assign io_ctl_r_rdata = 4'hf == addr[3:0] ? regs_15 : _GEN_17; // @[AXI4Lite2CTA.scala 79:{18,18}]
  assign io_ctl_r_rvalid = rvalid; // @[AXI4Lite2CTA.scala 90:19]
  assign io_ctl_r_rid = transaction_id; // @[AXI4Lite2CTA.scala 80:16]
  assign io_data_valid = input_valid & out_state; // @[AXI4Lite2CTA.scala 97:30]
  assign io_data_bits_host_wg_id = regs_1[4:0]; // @[AXI4Lite2CTA.scala 98:26]
  assign io_data_bits_host_num_wf = regs_2[2:0]; // @[AXI4Lite2CTA.scala 99:27]
  assign io_data_bits_host_wf_size = regs_3[9:0]; // @[AXI4Lite2CTA.scala 100:28]
  assign io_data_bits_host_start_pc = regs_4; // @[AXI4Lite2CTA.scala 101:29]
  assign io_data_bits_host_vgpr_size_total = regs_5[12:0]; // @[AXI4Lite2CTA.scala 102:36]
  assign io_data_bits_host_sgpr_size_total = regs_6[12:0]; // @[AXI4Lite2CTA.scala 103:36]
  assign io_data_bits_host_lds_size_total = regs_7[12:0]; // @[AXI4Lite2CTA.scala 104:35]
  assign io_data_bits_host_gds_size_total = regs_8[10:0]; // @[AXI4Lite2CTA.scala 105:35]
  assign io_data_bits_host_vgpr_size_per_wf = regs_9[12:0]; // @[AXI4Lite2CTA.scala 106:37]
  assign io_data_bits_host_sgpr_size_per_wf = regs_10[12:0]; // @[AXI4Lite2CTA.scala 107:37]
  assign io_rsp_ready = io_rsp_valid & ~regs_15[0]; // @[AXI4Lite2CTA.scala 53:20]
  always @(posedge clock) begin
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_0 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h0 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_0 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end else begin
        regs_0 <= _GEN_25;
      end
    end else begin
      regs_0 <= _GEN_25;
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_1 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h1 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_1 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_2 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h2 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_2 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_3 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h3 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_3 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_4 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h4 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_4 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_5 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h5 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_5 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_6 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h6 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_6 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_7 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h7 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_7 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_8 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h8 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_8 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_9 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'h9 == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_9 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_10 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'ha == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_10 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_11 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'hb == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_11 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_12 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'hc == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_12 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_13 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'hd == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_13 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_14 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'he == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_14 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end else begin
        regs_14 <= _GEN_2;
      end
    end else begin
      regs_14 <= _GEN_2;
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 50:21]
      regs_15 <= 32'h0; // @[AXI4Lite2CTA.scala 50:21]
    end else if (write) begin // @[AXI4Lite2CTA.scala 123:15]
      if (4'hf == addr[3:0]) begin // @[AXI4Lite2CTA.scala 124:16]
        regs_15 <= dataOut; // @[AXI4Lite2CTA.scala 124:16]
      end else begin
        regs_15 <= _GEN_1;
      end
    end else begin
      regs_15 <= _GEN_1;
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 60:22]
      state <= 3'h0; // @[AXI4Lite2CTA.scala 60:22]
    end else if (3'h0 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      if (io_ctl_aw_awvalid & _T_3) begin // @[AXI4Lite2CTA.scala 134:52]
        state <= 3'h3; // @[AXI4Lite2CTA.scala 135:15]
      end else if (io_ctl_ar_arvalid) begin // @[AXI4Lite2CTA.scala 137:36]
        state <= 3'h1; // @[AXI4Lite2CTA.scala 138:15]
      end
    end else if (3'h1 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      if (io_ctl_ar_arvalid & arready) begin // @[AXI4Lite2CTA.scala 145:41]
        state <= 3'h2; // @[AXI4Lite2CTA.scala 146:15]
      end
    end else if (3'h2 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      state <= _GEN_66;
    end else begin
      state <= _GEN_87;
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 62:24]
      awready <= 1'h0; // @[AXI4Lite2CTA.scala 62:24]
    end else if (!(3'h0 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (!(3'h1 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
        if (!(3'h2 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
          awready <= _GEN_85;
        end
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 63:23]
      wready <= 1'h0; // @[AXI4Lite2CTA.scala 63:23]
    end else if (!(3'h0 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (!(3'h1 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
        if (!(3'h2 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
          wready <= _GEN_88;
        end
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 64:23]
      bvalid <= 1'h0; // @[AXI4Lite2CTA.scala 64:23]
    end else if (3'h0 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      bvalid <= 1'h0; // @[AXI4Lite2CTA.scala 130:14]
    end else if (!(3'h1 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (!(3'h2 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
        bvalid <= _GEN_91;
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 67:24]
      arready <= 1'h0; // @[AXI4Lite2CTA.scala 67:24]
    end else if (!(3'h0 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (3'h1 == state) begin // @[AXI4Lite2CTA.scala 127:16]
        if (io_ctl_ar_arvalid & arready) begin // @[AXI4Lite2CTA.scala 145:41]
          arready <= 1'h0; // @[AXI4Lite2CTA.scala 149:17]
        end else begin
          arready <= 1'h1; // @[AXI4Lite2CTA.scala 144:15]
        end
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 68:23]
      rvalid <= 1'h0; // @[AXI4Lite2CTA.scala 68:23]
    end else if (3'h0 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      rvalid <= 1'h0; // @[AXI4Lite2CTA.scala 129:14]
    end else if (!(3'h1 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (3'h2 == state) begin // @[AXI4Lite2CTA.scala 127:16]
        rvalid <= _GEN_67;
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 71:21]
      addr <= 32'h0; // @[AXI4Lite2CTA.scala 71:21]
    end else if (!(3'h0 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (3'h1 == state) begin // @[AXI4Lite2CTA.scala 127:16]
        if (io_ctl_ar_arvalid & arready) begin // @[AXI4Lite2CTA.scala 145:41]
          addr <= {{2'd0}, io_ctl_ar_araddr[31:2]}; // @[AXI4Lite2CTA.scala 147:14]
        end
      end else if (!(3'h2 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
        addr <= _GEN_86;
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 74:22]
      write <= 1'h0; // @[AXI4Lite2CTA.scala 74:22]
    end else if (3'h0 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      write <= 1'h0; // @[AXI4Lite2CTA.scala 132:13]
    end else if (!(3'h1 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (!(3'h2 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
        write <= _GEN_90;
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 75:24]
      dataOut <= 32'h0; // @[AXI4Lite2CTA.scala 75:24]
    end else if (!(3'h0 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
      if (!(3'h1 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
        if (!(3'h2 == state)) begin // @[AXI4Lite2CTA.scala 127:16]
          dataOut <= _GEN_89;
        end
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 77:31]
      transaction_id <= 12'h0; // @[AXI4Lite2CTA.scala 77:31]
    end else if (3'h0 == state) begin // @[AXI4Lite2CTA.scala 127:16]
      if (io_ctl_aw_awvalid & _T_3) begin // @[AXI4Lite2CTA.scala 134:52]
        transaction_id <= io_ctl_aw_awid; // @[AXI4Lite2CTA.scala 136:24]
      end else if (io_ctl_ar_arvalid) begin // @[AXI4Lite2CTA.scala 137:36]
        transaction_id <= io_ctl_ar_arid; // @[AXI4Lite2CTA.scala 139:24]
      end else begin
        transaction_id <= 12'h0; // @[AXI4Lite2CTA.scala 133:22]
      end
    end
    if (reset) begin // @[AXI4Lite2CTA.scala 95:24]
      out_state <= 1'h0; // @[AXI4Lite2CTA.scala 95:24]
    end else if (~out_state) begin // @[AXI4Lite2CTA.scala 110:21]
      out_state <= _GEN_19;
    end else if (out_state) begin // @[AXI4Lite2CTA.scala 110:21]
      if (_T_5) begin // @[AXI4Lite2CTA.scala 117:26]
        out_state <= 1'h0; // @[AXI4Lite2CTA.scala 118:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  awready = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  wready = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  bvalid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  arready = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  rvalid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  addr = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  write = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  dataOut = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  transaction_id = _RAND_25[11:0];
  _RAND_26 = {1{`RANDOM}};
  out_state = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Adapter(
  input          clock,
  input          reset,
  input          io_AXI_master_bundle_aw_ready,
  output         io_AXI_master_bundle_aw_valid,
  output [3:0]   io_AXI_master_bundle_aw_bits_id,
  output [31:0]  io_AXI_master_bundle_aw_bits_addr,
  input          io_AXI_master_bundle_w_ready,
  output         io_AXI_master_bundle_w_valid,
  output [63:0]  io_AXI_master_bundle_w_bits_data,
  output [7:0]   io_AXI_master_bundle_w_bits_strb,
  output         io_AXI_master_bundle_w_bits_last,
  input          io_AXI_master_bundle_b_valid,
  input  [3:0]   io_AXI_master_bundle_b_bits_id,
  input          io_AXI_master_bundle_ar_ready,
  output         io_AXI_master_bundle_ar_valid,
  output [3:0]   io_AXI_master_bundle_ar_bits_id,
  output [31:0]  io_AXI_master_bundle_ar_bits_addr,
  output         io_AXI_master_bundle_r_ready,
  input          io_AXI_master_bundle_r_valid,
  input  [3:0]   io_AXI_master_bundle_r_bits_id,
  input  [63:0]  io_AXI_master_bundle_r_bits_data,
  input          io_AXI_master_bundle_r_bits_last,
  output         io_l2cache_outa_ready,
  input          io_l2cache_outa_valid,
  input  [2:0]   io_l2cache_outa_bits_opcode,
  input  [3:0]   io_l2cache_outa_bits_source,
  input  [31:0]  io_l2cache_outa_bits_address,
  input  [31:0]  io_l2cache_outa_bits_mask,
  input  [255:0] io_l2cache_outa_bits_data,
  input          io_l2cache_outd_ready,
  output         io_l2cache_outd_valid,
  output [2:0]   io_l2cache_outd_bits_opcode,
  output [3:0]   io_l2cache_outd_bits_source,
  output [255:0] io_l2cache_outd_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] counter_read; // @[AXI4Adapter.scala 42:27]
  reg [3:0] counter_write; // @[AXI4Adapter.scala 43:28]
  reg [3:0] buffer_read_0_id; // @[AXI4Adapter.scala 45:46]
  reg [63:0] buffer_read_0_data; // @[AXI4Adapter.scala 45:46]
  reg [3:0] buffer_read_1_id; // @[AXI4Adapter.scala 45:46]
  reg [63:0] buffer_read_1_data; // @[AXI4Adapter.scala 45:46]
  reg [3:0] buffer_read_2_id; // @[AXI4Adapter.scala 45:46]
  reg [63:0] buffer_read_2_data; // @[AXI4Adapter.scala 45:46]
  reg [3:0] buffer_read_3_id; // @[AXI4Adapter.scala 45:46]
  reg [63:0] buffer_read_3_data; // @[AXI4Adapter.scala 45:46]
  reg  buffer_read_valid; // @[AXI4Adapter.scala 46:32]
  reg  buffer_read_ready; // @[AXI4Adapter.scala 48:32]
  reg [7:0] buffer_write_0_mask; // @[AXI4Adapter.scala 49:46]
  reg [63:0] buffer_write_0_data; // @[AXI4Adapter.scala 49:46]
  reg [7:0] buffer_write_1_mask; // @[AXI4Adapter.scala 49:46]
  reg [63:0] buffer_write_1_data; // @[AXI4Adapter.scala 49:46]
  reg [7:0] buffer_write_2_mask; // @[AXI4Adapter.scala 49:46]
  reg [63:0] buffer_write_2_data; // @[AXI4Adapter.scala 49:46]
  reg [7:0] buffer_write_3_mask; // @[AXI4Adapter.scala 49:46]
  reg [63:0] buffer_write_3_data; // @[AXI4Adapter.scala 49:46]
  reg  buffer_write_valid; // @[AXI4Adapter.scala 50:33]
  wire  _io_AXI_master_bundle_aw_valid_T = io_l2cache_outa_bits_opcode == 3'h0; // @[AXI4Adapter.scala 55:65]
  wire  _io_AXI_master_bundle_aw_valid_T_1 = io_l2cache_outa_ready & io_l2cache_outa_valid; // @[Decoupled.scala 50:35]
  wire  _T = io_AXI_master_bundle_r_ready & io_AXI_master_bundle_r_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = buffer_read_valid & buffer_read_ready ? 1'h0 : buffer_read_valid; // @[AXI4Adapter.scala 91:53 92:22 46:32]
  wire  _GEN_1 = io_AXI_master_bundle_r_bits_last & _T | _GEN_0; // @[AXI4Adapter.scala 89:75 90:22]
  wire  buffer_read_busy = counter_read != 4'h0; // @[AXI4Adapter.scala 94:34]
  wire [3:0] _counter_read_T_1 = counter_read + 4'h1; // @[AXI4Adapter.scala 100:36]
  wire  _T_16 = io_AXI_master_bundle_aw_ready & io_AXI_master_bundle_aw_valid; // @[Decoupled.scala 50:35]
  wire  _T_18 = io_AXI_master_bundle_w_ready & io_AXI_master_bundle_w_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_20 = counter_write == 4'h3 & _T_18 ? 1'h0 : buffer_write_valid; // @[AXI4Adapter.scala 115:86 116:23 50:33]
  wire  _GEN_21 = _T_16 | _GEN_20; // @[AXI4Adapter.scala 113:38 114:24]
  reg  write_busy_reg; // @[AXI4Adapter.scala 118:29]
  wire  buffer_write_busy = write_busy_reg | counter_write != 4'h0 & counter_write != 4'h3; // @[AXI4Adapter.scala 119:37]
  wire [3:0] _counter_write_T_1 = counter_write + 4'h1; // @[AXI4Adapter.scala 124:38]
  wire [1:0] io_AXI_master_bundle_w_bits_data_truncIdx = counter_write[1:0]; // @[package.scala 31:49]
  wire [7:0] _io_AXI_master_bundle_w_bits_data_T_1_mask = io_AXI_master_bundle_w_bits_data_truncIdx == 2'h1 ?
    buffer_write_1_mask : buffer_write_0_mask; // @[package.scala 32:76]
  wire [63:0] _io_AXI_master_bundle_w_bits_data_T_1_data = io_AXI_master_bundle_w_bits_data_truncIdx == 2'h1 ?
    buffer_write_1_data : buffer_write_0_data; // @[package.scala 32:76]
  wire [7:0] _io_AXI_master_bundle_w_bits_data_T_3_mask = io_AXI_master_bundle_w_bits_data_truncIdx == 2'h2 ?
    buffer_write_2_mask : _io_AXI_master_bundle_w_bits_data_T_1_mask; // @[package.scala 32:76]
  wire [63:0] _io_AXI_master_bundle_w_bits_data_T_3_data = io_AXI_master_bundle_w_bits_data_truncIdx == 2'h2 ?
    buffer_write_2_data : _io_AXI_master_bundle_w_bits_data_T_1_data; // @[package.scala 32:76]
  wire [67:0] _io_l2cache_outd_bits_source_T = {buffer_read_0_id,buffer_read_0_data}; // @[AXI4Adapter.scala 150:120]
  wire  _io_l2cache_outd_bits_opcode_T = io_AXI_master_bundle_b_valid ? 1'h0 : 1'h1; // @[AXI4Adapter.scala 151:35]
  wire [67:0] _io_l2cache_outd_bits_data_T_3 = {buffer_read_1_id,buffer_read_1_data}; // @[AXI4Adapter.scala 152:93]
  wire [67:0] _io_l2cache_outd_bits_data_T_6 = {buffer_read_2_id,buffer_read_2_data}; // @[AXI4Adapter.scala 152:93]
  wire [67:0] _io_l2cache_outd_bits_data_T_9 = {buffer_read_3_id,buffer_read_3_data}; // @[AXI4Adapter.scala 152:93]
  wire [255:0] _io_l2cache_outd_bits_data_T_12 = {_io_l2cache_outd_bits_data_T_9[63:0],_io_l2cache_outd_bits_data_T_6[63
    :0],_io_l2cache_outd_bits_data_T_3[63:0],_io_l2cache_outd_bits_source_T[63:0]}; // @[Cat.scala 31:58]
  assign io_AXI_master_bundle_aw_valid = io_l2cache_outa_bits_opcode == 3'h0 & _io_AXI_master_bundle_aw_valid_T_1; // @[AXI4Adapter.scala 55:82]
  assign io_AXI_master_bundle_aw_bits_id = io_l2cache_outa_bits_source; // @[AXI4Adapter.scala 76:34]
  assign io_AXI_master_bundle_aw_bits_addr = io_l2cache_outa_bits_address; // @[AXI4Adapter.scala 72:37]
  assign io_AXI_master_bundle_w_valid = buffer_write_valid; // @[AXI4Adapter.scala 138:31]
  assign io_AXI_master_bundle_w_bits_data = io_AXI_master_bundle_w_bits_data_truncIdx == 2'h3 ? buffer_write_3_data :
    _io_AXI_master_bundle_w_bits_data_T_3_data; // @[package.scala 32:76]
  assign io_AXI_master_bundle_w_bits_strb = io_AXI_master_bundle_w_bits_data_truncIdx == 2'h3 ? buffer_write_3_mask :
    _io_AXI_master_bundle_w_bits_data_T_3_mask; // @[package.scala 32:76]
  assign io_AXI_master_bundle_w_bits_last = counter_write == 4'h3; // @[AXI4Adapter.scala 140:52]
  assign io_AXI_master_bundle_ar_valid = io_l2cache_outa_bits_opcode == 3'h4 & _io_AXI_master_bundle_aw_valid_T_1; // @[AXI4Adapter.scala 57:72]
  assign io_AXI_master_bundle_ar_bits_id = io_l2cache_outa_bits_source; // @[AXI4Adapter.scala 64:34]
  assign io_AXI_master_bundle_ar_bits_addr = io_l2cache_outa_bits_address; // @[AXI4Adapter.scala 59:37]
  assign io_AXI_master_bundle_r_ready = buffer_read_valid ? io_l2cache_outd_ready : 1'h1; // @[AXI4Adapter.scala 144:37]
  assign io_l2cache_outa_ready = ~buffer_write_busy & io_AXI_master_bundle_aw_ready & ~buffer_read_busy &
    io_AXI_master_bundle_ar_ready; // @[AXI4Adapter.scala 156:100]
  assign io_l2cache_outd_valid = io_AXI_master_bundle_b_valid | buffer_read_valid; // @[AXI4Adapter.scala 149:56]
  assign io_l2cache_outd_bits_opcode = {{2'd0}, _io_l2cache_outd_bits_opcode_T}; // @[AXI4Adapter.scala 151:30]
  assign io_l2cache_outd_bits_source = io_AXI_master_bundle_b_valid ? io_AXI_master_bundle_b_bits_id :
    _io_l2cache_outd_bits_source_T[67:64]; // @[AXI4Adapter.scala 150:36]
  assign io_l2cache_outd_bits_data = io_AXI_master_bundle_b_valid ? 256'h0 : _io_l2cache_outd_bits_data_T_12; // @[AXI4Adapter.scala 152:33]
  always @(posedge clock) begin
    if (reset) begin // @[AXI4Adapter.scala 42:27]
      counter_read <= 4'h0; // @[AXI4Adapter.scala 42:27]
    end else if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (io_AXI_master_bundle_r_bits_last) begin // @[AXI4Adapter.scala 97:43]
        counter_read <= 4'h0; // @[AXI4Adapter.scala 98:20]
      end else begin
        counter_read <= _counter_read_T_1; // @[AXI4Adapter.scala 100:20]
      end
    end
    if (reset) begin // @[AXI4Adapter.scala 43:28]
      counter_write <= 4'h0; // @[AXI4Adapter.scala 43:28]
    end else if (_T_18) begin // @[AXI4Adapter.scala 120:36]
      if (io_AXI_master_bundle_w_bits_last) begin // @[AXI4Adapter.scala 121:43]
        counter_write <= 4'h0; // @[AXI4Adapter.scala 122:21]
      end else begin
        counter_write <= _counter_write_T_1; // @[AXI4Adapter.scala 124:21]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h0 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_0_id <= io_AXI_master_bundle_r_bits_id; // @[AXI4Adapter.scala 106:29]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h0 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_0_data <= io_AXI_master_bundle_r_bits_data; // @[AXI4Adapter.scala 105:31]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h1 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_1_id <= io_AXI_master_bundle_r_bits_id; // @[AXI4Adapter.scala 106:29]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h1 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_1_data <= io_AXI_master_bundle_r_bits_data; // @[AXI4Adapter.scala 105:31]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h2 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_2_id <= io_AXI_master_bundle_r_bits_id; // @[AXI4Adapter.scala 106:29]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h2 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_2_data <= io_AXI_master_bundle_r_bits_data; // @[AXI4Adapter.scala 105:31]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h3 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_3_id <= io_AXI_master_bundle_r_bits_id; // @[AXI4Adapter.scala 106:29]
      end
    end
    if (_T) begin // @[AXI4Adapter.scala 96:36]
      if (_T & 4'h3 == counter_read) begin // @[AXI4Adapter.scala 104:74]
        buffer_read_3_data <= io_AXI_master_bundle_r_bits_data; // @[AXI4Adapter.scala 105:31]
      end
    end
    if (reset) begin // @[AXI4Adapter.scala 46:32]
      buffer_read_valid <= 1'h0; // @[AXI4Adapter.scala 46:32]
    end else begin
      buffer_read_valid <= _GEN_1;
    end
    buffer_read_ready <= reset | io_l2cache_outd_ready; // @[AXI4Adapter.scala 48:{32,32} 95:20]
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_0_mask <= io_l2cache_outa_bits_mask[7:0]; // @[AXI4Adapter.scala 132:16]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_0_data <= io_l2cache_outa_bits_data[63:0]; // @[AXI4Adapter.scala 130:15]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_1_mask <= io_l2cache_outa_bits_mask[15:8]; // @[AXI4Adapter.scala 132:16]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_1_data <= io_l2cache_outa_bits_data[127:64]; // @[AXI4Adapter.scala 130:15]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_2_mask <= io_l2cache_outa_bits_mask[23:16]; // @[AXI4Adapter.scala 132:16]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_2_data <= io_l2cache_outa_bits_data[191:128]; // @[AXI4Adapter.scala 130:15]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_3_mask <= io_l2cache_outa_bits_mask[31:24]; // @[AXI4Adapter.scala 132:16]
    end
    if (_io_AXI_master_bundle_aw_valid_T_1 & (_io_AXI_master_bundle_aw_valid_T | io_l2cache_outa_bits_opcode == 3'h1)
      ) begin // @[AXI4Adapter.scala 127:124]
      buffer_write_3_data <= io_l2cache_outa_bits_data[255:192]; // @[AXI4Adapter.scala 130:15]
    end
    if (reset) begin // @[AXI4Adapter.scala 50:33]
      buffer_write_valid <= 1'h0; // @[AXI4Adapter.scala 50:33]
    end else begin
      buffer_write_valid <= _GEN_21;
    end
    write_busy_reg <= io_AXI_master_bundle_aw_ready & io_AXI_master_bundle_aw_valid; // @[Decoupled.scala 50:35]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter_read = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  counter_write = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_read_0_id = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  buffer_read_0_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_read_1_id = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  buffer_read_1_data = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_read_2_id = _RAND_6[3:0];
  _RAND_7 = {2{`RANDOM}};
  buffer_read_2_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_read_3_id = _RAND_8[3:0];
  _RAND_9 = {2{`RANDOM}};
  buffer_read_3_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_read_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_read_ready = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_write_0_mask = _RAND_12[7:0];
  _RAND_13 = {2{`RANDOM}};
  buffer_write_0_data = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_write_1_mask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  buffer_write_1_data = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_write_2_mask = _RAND_16[7:0];
  _RAND_17 = {2{`RANDOM}};
  buffer_write_2_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_write_3_mask = _RAND_18[7:0];
  _RAND_19 = {2{`RANDOM}};
  buffer_write_3_data = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_write_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  write_busy_reg = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GPGPU_axi_top(
  input         clock,
  input         reset,
  input  [31:0] io_s_aw_awaddr,
  input  [2:0]  io_s_aw_awprot,
  input         io_s_aw_awvalid,
  output        io_s_aw_awready,
  input  [11:0] io_s_aw_awid,
  input  [31:0] io_s_w_wdata,
  input  [3:0]  io_s_w_wstrb,
  input         io_s_w_wvalid,
  output        io_s_w_wready,
  input  [11:0] io_s_w_wid,
  output [1:0]  io_s_b_bresp,
  output        io_s_b_bvalid,
  input         io_s_b_bready,
  output [11:0] io_s_b_bid,
  input  [31:0] io_s_ar_araddr,
  input  [2:0]  io_s_ar_arprot,
  input         io_s_ar_arvalid,
  output        io_s_ar_arready,
  input  [11:0] io_s_ar_arid,
  output [31:0] io_s_r_rdata,
  output [1:0]  io_s_r_rresp,
  output        io_s_r_rvalid,
  input         io_s_r_rready,
  output [11:0] io_s_r_rid,
  input         io_m_aw_ready,
  output        io_m_aw_valid,
  output [3:0]  io_m_aw_bits_id,
  output [31:0] io_m_aw_bits_addr,
  output [7:0]  io_m_aw_bits_len,
  output [2:0]  io_m_aw_bits_size,
  output [1:0]  io_m_aw_bits_burst,
  output        io_m_aw_bits_lock,
  output [3:0]  io_m_aw_bits_cache,
  output [2:0]  io_m_aw_bits_prot,
  output [3:0]  io_m_aw_bits_qos,
  input         io_m_w_ready,
  output        io_m_w_valid,
  output [63:0] io_m_w_bits_data,
  output [7:0]  io_m_w_bits_strb,
  output        io_m_w_bits_last,
  output        io_m_b_ready,
  input         io_m_b_valid,
  input  [3:0]  io_m_b_bits_id,
  input  [1:0]  io_m_b_bits_resp,
  input         io_m_ar_ready,
  output        io_m_ar_valid,
  output [3:0]  io_m_ar_bits_id,
  output [31:0] io_m_ar_bits_addr,
  output [7:0]  io_m_ar_bits_len,
  output [2:0]  io_m_ar_bits_size,
  output [1:0]  io_m_ar_bits_burst,
  output        io_m_ar_bits_lock,
  output [3:0]  io_m_ar_bits_cache,
  output [2:0]  io_m_ar_bits_prot,
  output [3:0]  io_m_ar_bits_qos,
  output        io_m_r_ready,
  input         io_m_r_valid,
  input  [3:0]  io_m_r_bits_id,
  input  [63:0] io_m_r_bits_data,
  input  [1:0]  io_m_r_bits_resp,
  input         io_m_r_bits_last
);
  wire  gpgpu_top_clock; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_reset; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_host_req_ready; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_host_req_valid; // @[GPGPU_top.scala 99:23]
  wire [4:0] gpgpu_top_io_host_req_bits_host_wg_id; // @[GPGPU_top.scala 99:23]
  wire [2:0] gpgpu_top_io_host_req_bits_host_num_wf; // @[GPGPU_top.scala 99:23]
  wire [9:0] gpgpu_top_io_host_req_bits_host_wf_size; // @[GPGPU_top.scala 99:23]
  wire [31:0] gpgpu_top_io_host_req_bits_host_start_pc; // @[GPGPU_top.scala 99:23]
  wire [12:0] gpgpu_top_io_host_req_bits_host_vgpr_size_total; // @[GPGPU_top.scala 99:23]
  wire [12:0] gpgpu_top_io_host_req_bits_host_sgpr_size_total; // @[GPGPU_top.scala 99:23]
  wire [12:0] gpgpu_top_io_host_req_bits_host_lds_size_total; // @[GPGPU_top.scala 99:23]
  wire [10:0] gpgpu_top_io_host_req_bits_host_gds_size_total; // @[GPGPU_top.scala 99:23]
  wire [12:0] gpgpu_top_io_host_req_bits_host_vgpr_size_per_wf; // @[GPGPU_top.scala 99:23]
  wire [12:0] gpgpu_top_io_host_req_bits_host_sgpr_size_per_wf; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_host_rsp_ready; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_host_rsp_valid; // @[GPGPU_top.scala 99:23]
  wire [4:0] gpgpu_top_io_host_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_out_a_ready; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_out_a_valid; // @[GPGPU_top.scala 99:23]
  wire [2:0] gpgpu_top_io_out_a_bits_opcode; // @[GPGPU_top.scala 99:23]
  wire [3:0] gpgpu_top_io_out_a_bits_source; // @[GPGPU_top.scala 99:23]
  wire [31:0] gpgpu_top_io_out_a_bits_address; // @[GPGPU_top.scala 99:23]
  wire [31:0] gpgpu_top_io_out_a_bits_mask; // @[GPGPU_top.scala 99:23]
  wire [255:0] gpgpu_top_io_out_a_bits_data; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_out_d_ready; // @[GPGPU_top.scala 99:23]
  wire  gpgpu_top_io_out_d_valid; // @[GPGPU_top.scala 99:23]
  wire [2:0] gpgpu_top_io_out_d_bits_opcode; // @[GPGPU_top.scala 99:23]
  wire [3:0] gpgpu_top_io_out_d_bits_source; // @[GPGPU_top.scala 99:23]
  wire [255:0] gpgpu_top_io_out_d_bits_data; // @[GPGPU_top.scala 99:23]
  wire  axi_lite_adapter_clock; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_reset; // @[GPGPU_top.scala 100:30]
  wire [31:0] axi_lite_adapter_io_ctl_aw_awaddr; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_aw_awvalid; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_aw_awready; // @[GPGPU_top.scala 100:30]
  wire [11:0] axi_lite_adapter_io_ctl_aw_awid; // @[GPGPU_top.scala 100:30]
  wire [31:0] axi_lite_adapter_io_ctl_w_wdata; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_w_wvalid; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_w_wready; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_b_bvalid; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_b_bready; // @[GPGPU_top.scala 100:30]
  wire [11:0] axi_lite_adapter_io_ctl_b_bid; // @[GPGPU_top.scala 100:30]
  wire [31:0] axi_lite_adapter_io_ctl_ar_araddr; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_ar_arvalid; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_ar_arready; // @[GPGPU_top.scala 100:30]
  wire [11:0] axi_lite_adapter_io_ctl_ar_arid; // @[GPGPU_top.scala 100:30]
  wire [31:0] axi_lite_adapter_io_ctl_r_rdata; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_r_rvalid; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_ctl_r_rready; // @[GPGPU_top.scala 100:30]
  wire [11:0] axi_lite_adapter_io_ctl_r_rid; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_data_ready; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_data_valid; // @[GPGPU_top.scala 100:30]
  wire [4:0] axi_lite_adapter_io_data_bits_host_wg_id; // @[GPGPU_top.scala 100:30]
  wire [2:0] axi_lite_adapter_io_data_bits_host_num_wf; // @[GPGPU_top.scala 100:30]
  wire [9:0] axi_lite_adapter_io_data_bits_host_wf_size; // @[GPGPU_top.scala 100:30]
  wire [31:0] axi_lite_adapter_io_data_bits_host_start_pc; // @[GPGPU_top.scala 100:30]
  wire [12:0] axi_lite_adapter_io_data_bits_host_vgpr_size_total; // @[GPGPU_top.scala 100:30]
  wire [12:0] axi_lite_adapter_io_data_bits_host_sgpr_size_total; // @[GPGPU_top.scala 100:30]
  wire [12:0] axi_lite_adapter_io_data_bits_host_lds_size_total; // @[GPGPU_top.scala 100:30]
  wire [10:0] axi_lite_adapter_io_data_bits_host_gds_size_total; // @[GPGPU_top.scala 100:30]
  wire [12:0] axi_lite_adapter_io_data_bits_host_vgpr_size_per_wf; // @[GPGPU_top.scala 100:30]
  wire [12:0] axi_lite_adapter_io_data_bits_host_sgpr_size_per_wf; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_rsp_ready; // @[GPGPU_top.scala 100:30]
  wire  axi_lite_adapter_io_rsp_valid; // @[GPGPU_top.scala 100:30]
  wire [4:0] axi_lite_adapter_io_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 100:30]
  wire  axi_adapter_clock; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_reset; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_aw_ready; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_aw_valid; // @[GPGPU_top.scala 101:25]
  wire [3:0] axi_adapter_io_AXI_master_bundle_aw_bits_id; // @[GPGPU_top.scala 101:25]
  wire [31:0] axi_adapter_io_AXI_master_bundle_aw_bits_addr; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_w_ready; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_w_valid; // @[GPGPU_top.scala 101:25]
  wire [63:0] axi_adapter_io_AXI_master_bundle_w_bits_data; // @[GPGPU_top.scala 101:25]
  wire [7:0] axi_adapter_io_AXI_master_bundle_w_bits_strb; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_w_bits_last; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_b_valid; // @[GPGPU_top.scala 101:25]
  wire [3:0] axi_adapter_io_AXI_master_bundle_b_bits_id; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_ar_ready; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_ar_valid; // @[GPGPU_top.scala 101:25]
  wire [3:0] axi_adapter_io_AXI_master_bundle_ar_bits_id; // @[GPGPU_top.scala 101:25]
  wire [31:0] axi_adapter_io_AXI_master_bundle_ar_bits_addr; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_r_ready; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_r_valid; // @[GPGPU_top.scala 101:25]
  wire [3:0] axi_adapter_io_AXI_master_bundle_r_bits_id; // @[GPGPU_top.scala 101:25]
  wire [63:0] axi_adapter_io_AXI_master_bundle_r_bits_data; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_AXI_master_bundle_r_bits_last; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_l2cache_outa_ready; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_l2cache_outa_valid; // @[GPGPU_top.scala 101:25]
  wire [2:0] axi_adapter_io_l2cache_outa_bits_opcode; // @[GPGPU_top.scala 101:25]
  wire [3:0] axi_adapter_io_l2cache_outa_bits_source; // @[GPGPU_top.scala 101:25]
  wire [31:0] axi_adapter_io_l2cache_outa_bits_address; // @[GPGPU_top.scala 101:25]
  wire [31:0] axi_adapter_io_l2cache_outa_bits_mask; // @[GPGPU_top.scala 101:25]
  wire [255:0] axi_adapter_io_l2cache_outa_bits_data; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_l2cache_outd_ready; // @[GPGPU_top.scala 101:25]
  wire  axi_adapter_io_l2cache_outd_valid; // @[GPGPU_top.scala 101:25]
  wire [2:0] axi_adapter_io_l2cache_outd_bits_opcode; // @[GPGPU_top.scala 101:25]
  wire [3:0] axi_adapter_io_l2cache_outd_bits_source; // @[GPGPU_top.scala 101:25]
  wire [255:0] axi_adapter_io_l2cache_outd_bits_data; // @[GPGPU_top.scala 101:25]
  GPGPU_top gpgpu_top ( // @[GPGPU_top.scala 99:23]
    .clock(gpgpu_top_clock),
    .reset(gpgpu_top_reset),
    .io_host_req_ready(gpgpu_top_io_host_req_ready),
    .io_host_req_valid(gpgpu_top_io_host_req_valid),
    .io_host_req_bits_host_wg_id(gpgpu_top_io_host_req_bits_host_wg_id),
    .io_host_req_bits_host_num_wf(gpgpu_top_io_host_req_bits_host_num_wf),
    .io_host_req_bits_host_wf_size(gpgpu_top_io_host_req_bits_host_wf_size),
    .io_host_req_bits_host_start_pc(gpgpu_top_io_host_req_bits_host_start_pc),
    .io_host_req_bits_host_vgpr_size_total(gpgpu_top_io_host_req_bits_host_vgpr_size_total),
    .io_host_req_bits_host_sgpr_size_total(gpgpu_top_io_host_req_bits_host_sgpr_size_total),
    .io_host_req_bits_host_lds_size_total(gpgpu_top_io_host_req_bits_host_lds_size_total),
    .io_host_req_bits_host_gds_size_total(gpgpu_top_io_host_req_bits_host_gds_size_total),
    .io_host_req_bits_host_vgpr_size_per_wf(gpgpu_top_io_host_req_bits_host_vgpr_size_per_wf),
    .io_host_req_bits_host_sgpr_size_per_wf(gpgpu_top_io_host_req_bits_host_sgpr_size_per_wf),
    .io_host_rsp_ready(gpgpu_top_io_host_rsp_ready),
    .io_host_rsp_valid(gpgpu_top_io_host_rsp_valid),
    .io_host_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id(
      gpgpu_top_io_host_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id),
    .io_out_a_ready(gpgpu_top_io_out_a_ready),
    .io_out_a_valid(gpgpu_top_io_out_a_valid),
    .io_out_a_bits_opcode(gpgpu_top_io_out_a_bits_opcode),
    .io_out_a_bits_source(gpgpu_top_io_out_a_bits_source),
    .io_out_a_bits_address(gpgpu_top_io_out_a_bits_address),
    .io_out_a_bits_mask(gpgpu_top_io_out_a_bits_mask),
    .io_out_a_bits_data(gpgpu_top_io_out_a_bits_data),
    .io_out_d_ready(gpgpu_top_io_out_d_ready),
    .io_out_d_valid(gpgpu_top_io_out_d_valid),
    .io_out_d_bits_opcode(gpgpu_top_io_out_d_bits_opcode),
    .io_out_d_bits_source(gpgpu_top_io_out_d_bits_source),
    .io_out_d_bits_data(gpgpu_top_io_out_d_bits_data)
  );
  AXI4Lite2CTA axi_lite_adapter ( // @[GPGPU_top.scala 100:30]
    .clock(axi_lite_adapter_clock),
    .reset(axi_lite_adapter_reset),
    .io_ctl_aw_awaddr(axi_lite_adapter_io_ctl_aw_awaddr),
    .io_ctl_aw_awvalid(axi_lite_adapter_io_ctl_aw_awvalid),
    .io_ctl_aw_awready(axi_lite_adapter_io_ctl_aw_awready),
    .io_ctl_aw_awid(axi_lite_adapter_io_ctl_aw_awid),
    .io_ctl_w_wdata(axi_lite_adapter_io_ctl_w_wdata),
    .io_ctl_w_wvalid(axi_lite_adapter_io_ctl_w_wvalid),
    .io_ctl_w_wready(axi_lite_adapter_io_ctl_w_wready),
    .io_ctl_b_bvalid(axi_lite_adapter_io_ctl_b_bvalid),
    .io_ctl_b_bready(axi_lite_adapter_io_ctl_b_bready),
    .io_ctl_b_bid(axi_lite_adapter_io_ctl_b_bid),
    .io_ctl_ar_araddr(axi_lite_adapter_io_ctl_ar_araddr),
    .io_ctl_ar_arvalid(axi_lite_adapter_io_ctl_ar_arvalid),
    .io_ctl_ar_arready(axi_lite_adapter_io_ctl_ar_arready),
    .io_ctl_ar_arid(axi_lite_adapter_io_ctl_ar_arid),
    .io_ctl_r_rdata(axi_lite_adapter_io_ctl_r_rdata),
    .io_ctl_r_rvalid(axi_lite_adapter_io_ctl_r_rvalid),
    .io_ctl_r_rready(axi_lite_adapter_io_ctl_r_rready),
    .io_ctl_r_rid(axi_lite_adapter_io_ctl_r_rid),
    .io_data_ready(axi_lite_adapter_io_data_ready),
    .io_data_valid(axi_lite_adapter_io_data_valid),
    .io_data_bits_host_wg_id(axi_lite_adapter_io_data_bits_host_wg_id),
    .io_data_bits_host_num_wf(axi_lite_adapter_io_data_bits_host_num_wf),
    .io_data_bits_host_wf_size(axi_lite_adapter_io_data_bits_host_wf_size),
    .io_data_bits_host_start_pc(axi_lite_adapter_io_data_bits_host_start_pc),
    .io_data_bits_host_vgpr_size_total(axi_lite_adapter_io_data_bits_host_vgpr_size_total),
    .io_data_bits_host_sgpr_size_total(axi_lite_adapter_io_data_bits_host_sgpr_size_total),
    .io_data_bits_host_lds_size_total(axi_lite_adapter_io_data_bits_host_lds_size_total),
    .io_data_bits_host_gds_size_total(axi_lite_adapter_io_data_bits_host_gds_size_total),
    .io_data_bits_host_vgpr_size_per_wf(axi_lite_adapter_io_data_bits_host_vgpr_size_per_wf),
    .io_data_bits_host_sgpr_size_per_wf(axi_lite_adapter_io_data_bits_host_sgpr_size_per_wf),
    .io_rsp_ready(axi_lite_adapter_io_rsp_ready),
    .io_rsp_valid(axi_lite_adapter_io_rsp_valid),
    .io_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id(
      axi_lite_adapter_io_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id)
  );
  AXI4Adapter axi_adapter ( // @[GPGPU_top.scala 101:25]
    .clock(axi_adapter_clock),
    .reset(axi_adapter_reset),
    .io_AXI_master_bundle_aw_ready(axi_adapter_io_AXI_master_bundle_aw_ready),
    .io_AXI_master_bundle_aw_valid(axi_adapter_io_AXI_master_bundle_aw_valid),
    .io_AXI_master_bundle_aw_bits_id(axi_adapter_io_AXI_master_bundle_aw_bits_id),
    .io_AXI_master_bundle_aw_bits_addr(axi_adapter_io_AXI_master_bundle_aw_bits_addr),
    .io_AXI_master_bundle_w_ready(axi_adapter_io_AXI_master_bundle_w_ready),
    .io_AXI_master_bundle_w_valid(axi_adapter_io_AXI_master_bundle_w_valid),
    .io_AXI_master_bundle_w_bits_data(axi_adapter_io_AXI_master_bundle_w_bits_data),
    .io_AXI_master_bundle_w_bits_strb(axi_adapter_io_AXI_master_bundle_w_bits_strb),
    .io_AXI_master_bundle_w_bits_last(axi_adapter_io_AXI_master_bundle_w_bits_last),
    .io_AXI_master_bundle_b_valid(axi_adapter_io_AXI_master_bundle_b_valid),
    .io_AXI_master_bundle_b_bits_id(axi_adapter_io_AXI_master_bundle_b_bits_id),
    .io_AXI_master_bundle_ar_ready(axi_adapter_io_AXI_master_bundle_ar_ready),
    .io_AXI_master_bundle_ar_valid(axi_adapter_io_AXI_master_bundle_ar_valid),
    .io_AXI_master_bundle_ar_bits_id(axi_adapter_io_AXI_master_bundle_ar_bits_id),
    .io_AXI_master_bundle_ar_bits_addr(axi_adapter_io_AXI_master_bundle_ar_bits_addr),
    .io_AXI_master_bundle_r_ready(axi_adapter_io_AXI_master_bundle_r_ready),
    .io_AXI_master_bundle_r_valid(axi_adapter_io_AXI_master_bundle_r_valid),
    .io_AXI_master_bundle_r_bits_id(axi_adapter_io_AXI_master_bundle_r_bits_id),
    .io_AXI_master_bundle_r_bits_data(axi_adapter_io_AXI_master_bundle_r_bits_data),
    .io_AXI_master_bundle_r_bits_last(axi_adapter_io_AXI_master_bundle_r_bits_last),
    .io_l2cache_outa_ready(axi_adapter_io_l2cache_outa_ready),
    .io_l2cache_outa_valid(axi_adapter_io_l2cache_outa_valid),
    .io_l2cache_outa_bits_opcode(axi_adapter_io_l2cache_outa_bits_opcode),
    .io_l2cache_outa_bits_source(axi_adapter_io_l2cache_outa_bits_source),
    .io_l2cache_outa_bits_address(axi_adapter_io_l2cache_outa_bits_address),
    .io_l2cache_outa_bits_mask(axi_adapter_io_l2cache_outa_bits_mask),
    .io_l2cache_outa_bits_data(axi_adapter_io_l2cache_outa_bits_data),
    .io_l2cache_outd_ready(axi_adapter_io_l2cache_outd_ready),
    .io_l2cache_outd_valid(axi_adapter_io_l2cache_outd_valid),
    .io_l2cache_outd_bits_opcode(axi_adapter_io_l2cache_outd_bits_opcode),
    .io_l2cache_outd_bits_source(axi_adapter_io_l2cache_outd_bits_source),
    .io_l2cache_outd_bits_data(axi_adapter_io_l2cache_outd_bits_data)
  );
  assign io_s_aw_awready = axi_lite_adapter_io_ctl_aw_awready; // @[GPGPU_top.scala 102:26]
  assign io_s_w_wready = axi_lite_adapter_io_ctl_w_wready; // @[GPGPU_top.scala 102:26]
  assign io_s_b_bresp = 2'h0; // @[GPGPU_top.scala 102:26]
  assign io_s_b_bvalid = axi_lite_adapter_io_ctl_b_bvalid; // @[GPGPU_top.scala 102:26]
  assign io_s_b_bid = axi_lite_adapter_io_ctl_b_bid; // @[GPGPU_top.scala 102:26]
  assign io_s_ar_arready = axi_lite_adapter_io_ctl_ar_arready; // @[GPGPU_top.scala 102:26]
  assign io_s_r_rdata = axi_lite_adapter_io_ctl_r_rdata; // @[GPGPU_top.scala 102:26]
  assign io_s_r_rresp = 2'h0; // @[GPGPU_top.scala 102:26]
  assign io_s_r_rvalid = axi_lite_adapter_io_ctl_r_rvalid; // @[GPGPU_top.scala 102:26]
  assign io_s_r_rid = axi_lite_adapter_io_ctl_r_rid; // @[GPGPU_top.scala 102:26]
  assign io_m_aw_valid = axi_adapter_io_AXI_master_bundle_aw_valid; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_id = axi_adapter_io_AXI_master_bundle_aw_bits_id; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_addr = axi_adapter_io_AXI_master_bundle_aw_bits_addr; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_len = 8'h3; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_size = 3'h3; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_burst = 2'h1; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_lock = 1'h0; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_cache = 4'h6; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_prot = 3'h0; // @[GPGPU_top.scala 103:35]
  assign io_m_aw_bits_qos = 4'h0; // @[GPGPU_top.scala 103:35]
  assign io_m_w_valid = axi_adapter_io_AXI_master_bundle_w_valid; // @[GPGPU_top.scala 103:35]
  assign io_m_w_bits_data = axi_adapter_io_AXI_master_bundle_w_bits_data; // @[GPGPU_top.scala 103:35]
  assign io_m_w_bits_strb = axi_adapter_io_AXI_master_bundle_w_bits_strb; // @[GPGPU_top.scala 103:35]
  assign io_m_w_bits_last = axi_adapter_io_AXI_master_bundle_w_bits_last; // @[GPGPU_top.scala 103:35]
  assign io_m_b_ready = 1'h1; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_valid = axi_adapter_io_AXI_master_bundle_ar_valid; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_id = axi_adapter_io_AXI_master_bundle_ar_bits_id; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_addr = axi_adapter_io_AXI_master_bundle_ar_bits_addr; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_len = 8'h3; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_size = 3'h3; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_burst = 2'h1; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_lock = 1'h0; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_cache = 4'h6; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_prot = 3'h0; // @[GPGPU_top.scala 103:35]
  assign io_m_ar_bits_qos = 4'h0; // @[GPGPU_top.scala 103:35]
  assign io_m_r_ready = axi_adapter_io_AXI_master_bundle_r_ready; // @[GPGPU_top.scala 103:35]
  assign gpgpu_top_clock = clock;
  assign gpgpu_top_reset = reset;
  assign gpgpu_top_io_host_req_valid = axi_lite_adapter_io_data_valid; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_wg_id = axi_lite_adapter_io_data_bits_host_wg_id; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_num_wf = axi_lite_adapter_io_data_bits_host_num_wf; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_wf_size = axi_lite_adapter_io_data_bits_host_wf_size; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_start_pc = axi_lite_adapter_io_data_bits_host_start_pc; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_vgpr_size_total = axi_lite_adapter_io_data_bits_host_vgpr_size_total; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_sgpr_size_total = axi_lite_adapter_io_data_bits_host_sgpr_size_total; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_lds_size_total = axi_lite_adapter_io_data_bits_host_lds_size_total; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_gds_size_total = axi_lite_adapter_io_data_bits_host_gds_size_total; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_vgpr_size_per_wf = axi_lite_adapter_io_data_bits_host_vgpr_size_per_wf; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_req_bits_host_sgpr_size_per_wf = axi_lite_adapter_io_data_bits_host_sgpr_size_per_wf; // @[GPGPU_top.scala 106:24]
  assign gpgpu_top_io_host_rsp_ready = axi_lite_adapter_io_rsp_ready; // @[GPGPU_top.scala 107:24]
  assign gpgpu_top_io_out_a_ready = axi_adapter_io_l2cache_outa_ready; // @[GPGPU_top.scala 104:21]
  assign gpgpu_top_io_out_d_valid = axi_adapter_io_l2cache_outd_valid; // @[GPGPU_top.scala 105:21]
  assign gpgpu_top_io_out_d_bits_opcode = axi_adapter_io_l2cache_outd_bits_opcode; // @[GPGPU_top.scala 105:21]
  assign gpgpu_top_io_out_d_bits_source = axi_adapter_io_l2cache_outd_bits_source; // @[GPGPU_top.scala 105:21]
  assign gpgpu_top_io_out_d_bits_data = axi_adapter_io_l2cache_outd_bits_data; // @[GPGPU_top.scala 105:21]
  assign axi_lite_adapter_clock = clock;
  assign axi_lite_adapter_reset = reset;
  assign axi_lite_adapter_io_ctl_aw_awaddr = io_s_aw_awaddr; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_aw_awvalid = io_s_aw_awvalid; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_aw_awid = io_s_aw_awid; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_w_wdata = io_s_w_wdata; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_w_wvalid = io_s_w_wvalid; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_b_bready = io_s_b_bready; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_ar_araddr = io_s_ar_araddr; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_ar_arvalid = io_s_ar_arvalid; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_ar_arid = io_s_ar_arid; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_ctl_r_rready = io_s_r_rready; // @[GPGPU_top.scala 102:26]
  assign axi_lite_adapter_io_data_ready = gpgpu_top_io_host_req_ready; // @[GPGPU_top.scala 106:24]
  assign axi_lite_adapter_io_rsp_valid = gpgpu_top_io_host_rsp_valid; // @[GPGPU_top.scala 107:24]
  assign axi_lite_adapter_io_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id =
    gpgpu_top_io_host_rsp_bits_inflight_wg_buffer_host_wf_done_wg_id; // @[GPGPU_top.scala 107:24]
  assign axi_adapter_clock = clock;
  assign axi_adapter_reset = reset;
  assign axi_adapter_io_AXI_master_bundle_aw_ready = io_m_aw_ready; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_w_ready = io_m_w_ready; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_b_valid = io_m_b_valid; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_b_bits_id = io_m_b_bits_id; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_ar_ready = io_m_ar_ready; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_r_valid = io_m_r_valid; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_r_bits_id = io_m_r_bits_id; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_r_bits_data = io_m_r_bits_data; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_AXI_master_bundle_r_bits_last = io_m_r_bits_last; // @[GPGPU_top.scala 103:35]
  assign axi_adapter_io_l2cache_outa_valid = gpgpu_top_io_out_a_valid; // @[GPGPU_top.scala 104:21]
  assign axi_adapter_io_l2cache_outa_bits_opcode = gpgpu_top_io_out_a_bits_opcode; // @[GPGPU_top.scala 104:21]
  assign axi_adapter_io_l2cache_outa_bits_source = gpgpu_top_io_out_a_bits_source; // @[GPGPU_top.scala 104:21]
  assign axi_adapter_io_l2cache_outa_bits_address = gpgpu_top_io_out_a_bits_address; // @[GPGPU_top.scala 104:21]
  assign axi_adapter_io_l2cache_outa_bits_mask = gpgpu_top_io_out_a_bits_mask; // @[GPGPU_top.scala 104:21]
  assign axi_adapter_io_l2cache_outa_bits_data = gpgpu_top_io_out_a_bits_data; // @[GPGPU_top.scala 104:21]
  assign axi_adapter_io_l2cache_outd_ready = gpgpu_top_io_out_d_ready; // @[GPGPU_top.scala 105:21]
endmodule
